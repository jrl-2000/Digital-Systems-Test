module Fictitious_CPU(Input, Output);

	input [7:0] Input;
	output [15:0] Output;
	
	// Fictitious CPU

endmodule