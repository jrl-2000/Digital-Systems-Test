
//Verilog file of module Circuit298


`timescale 1 ns / 1ns

module s298_unfolded(Clock,
reset,
g0,
g1,
g2,
g117,
g132,
g66,
g118,
g133,
g67,
Circuit298_wire_3,
Circuit298_wire_5,
Circuit298_wire_7,
Circuit298_wire_9,
Circuit298_wire_11,
Circuit298_wire_13,
Circuit298_wire_15,
Circuit298_wire_17,
Circuit298_wire_19,
Circuit298_wire_21,
Circuit298_wire_23,
Circuit298_wire_26,
Circuit298_wire_28,
Circuit298_wire_30,
Circuit298_wire_32,
Circuit298_wire_34,
Circuit298_wire_36,
Circuit298_wire_38,
Circuit298_wire_40,
Circuit298_wire_42,
Circuit298_wire_44,
Circuit298_wire_46,
Circuit298_wire_48,
Circuit298_wire_50,
Circuit298_wire_52,
/////////////////////
Circuit298_wire_2_out,
Circuit298_wire_4_out,
Circuit298_wire_6_out,
Circuit298_wire_8_out,
Circuit298_wire_10_out,
Circuit298_wire_12_out,
Circuit298_wire_14_out,
Circuit298_wire_16_out,
Circuit298_wire_18_out,
Circuit298_wire_20_out,
Circuit298_wire_22_out,
Circuit298_wire_25_out,
Circuit298_wire_27_out,
Circuit298_wire_29_out,
Circuit298_wire_31_out,
Circuit298_wire_33_out,
Circuit298_wire_35_out,
Circuit298_wire_37_out,
Circuit298_wire_39_out,
Circuit298_wire_41_out,
Circuit298_wire_43_out,
Circuit298_wire_45_out,
Circuit298_wire_47_out,
Circuit298_wire_49_out,
Circuit298_wire_51_out
);
  input  Clock;
  input  reset;
  input  g0;
  input  g1;
  input  g2;
  input  Circuit298_wire_3; 
  input  Circuit298_wire_5; 
  input  Circuit298_wire_7; 
  input  Circuit298_wire_9; 
  input  Circuit298_wire_11;
  input  Circuit298_wire_13;
  input  Circuit298_wire_15;
  input  Circuit298_wire_17;
  input  Circuit298_wire_19;
  input  Circuit298_wire_21;
  input  Circuit298_wire_23;
  input  Circuit298_wire_26;
  input  Circuit298_wire_28;
  input  Circuit298_wire_30;
  input  Circuit298_wire_32;
  input  Circuit298_wire_34;
  input  Circuit298_wire_36;
  input  Circuit298_wire_38;
  input  Circuit298_wire_40;
  input  Circuit298_wire_42;
  input  Circuit298_wire_44;
  input  Circuit298_wire_46;
  input  Circuit298_wire_48;
  input  Circuit298_wire_50;
  input  Circuit298_wire_52;

  
  
  output Circuit298_wire_2_out;
  output Circuit298_wire_4_out; 
  output Circuit298_wire_6_out;
  output Circuit298_wire_8_out; 
  output Circuit298_wire_10_out;
  output Circuit298_wire_12_out;
  output Circuit298_wire_14_out;
  output Circuit298_wire_16_out;
  output Circuit298_wire_18_out;
  output Circuit298_wire_20_out;
  output Circuit298_wire_22_out;
  output Circuit298_wire_25_out;
  output Circuit298_wire_27_out;
  output Circuit298_wire_29_out;
  output Circuit298_wire_31_out;
  output Circuit298_wire_33_out;
  output Circuit298_wire_35_out;
  output Circuit298_wire_37_out;
  output Circuit298_wire_39_out;
  output Circuit298_wire_41_out;
  output Circuit298_wire_43_out;
  output Circuit298_wire_45_out;
  output Circuit298_wire_47_out;
  output Circuit298_wire_49_out;
  output Circuit298_wire_51_out;
  output g117;
  output g132;
  output g66;
  output g118;
  output g133;
  output g67;

wire
Circuit298_wire_1,
//Circuit298_wire_2,
//Circuit298_wire_3,
//Circuit298_wire_4,
//Circuit298_wire_5,
//Circuit298_wire_6,
//Circuit298_wire_7,
//Circuit298_wire_8,
//Circuit298_wire_9,
//Circuit298_wire_10,
//Circuit298_wire_11,
//Circuit298_wire_12,
//Circuit298_wire_13,
//Circuit298_wire_14,
//Circuit298_wire_15,
//Circuit298_wire_16,
//Circuit298_wire_17,
//Circuit298_wire_18,
//Circuit298_wire_19,
//Circuit298_wire_20,
//Circuit298_wire_21,
//Circuit298_wire_22,
//Circuit298_wire_23,
Circuit298_wire_24,
//Circuit298_wire_25,
//Circuit298_wire_26,
//Circuit298_wire_27,
//Circuit298_wire_28,
//Circuit298_wire_29,
//Circuit298_wire_30,
//Circuit298_wire_31,
//Circuit298_wire_32,
//Circuit298_wire_33,
//Circuit298_wire_34,
//Circuit298_wire_35,
//Circuit298_wire_36,
//Circuit298_wire_37,
//Circuit298_wire_38,
//Circuit298_wire_39,
//Circuit298_wire_40,
//Circuit298_wire_41,
//Circuit298_wire_42,
//Circuit298_wire_43,
//Circuit298_wire_44,
//Circuit298_wire_45,
//Circuit298_wire_46,
//Circuit298_wire_47,
//Circuit298_wire_48,
//Circuit298_wire_49,
//Circuit298_wire_50,
//Circuit298_wire_51,
//Circuit298_wire_52,
Circuit298_wire_53,
Circuit298_wire_54,
Circuit298_wire_55,
Circuit298_wire_56,
Circuit298_wire_57,
Circuit298_wire_58,
Circuit298_wire_59,
Circuit298_wire_60,
Circuit298_wire_61,
Circuit298_wire_62,
Circuit298_wire_63,
Circuit298_wire_64,
Circuit298_wire_65,
Circuit298_wire_66,
Circuit298_wire_67,
Circuit298_wire_68,
Circuit298_wire_69,
Circuit298_wire_70,
Circuit298_wire_71,
Circuit298_wire_72,
Circuit298_wire_73,
Circuit298_wire_74,
Circuit298_wire_75,
Circuit298_wire_76,
Circuit298_wire_77,
Circuit298_wire_78,
Circuit298_wire_79,
Circuit298_wire_80,
Circuit298_wire_81,
Circuit298_wire_82,
Circuit298_wire_83,
Circuit298_wire_84,
Circuit298_wire_85,
Circuit298_wire_86,
Circuit298_wire_87,
Circuit298_wire_88,
Circuit298_wire_89,
Circuit298_wire_90,
Circuit298_wire_91,
Circuit298_wire_92,
Circuit298_wire_93,
Circuit298_wire_94,
Circuit298_wire_95,
Circuit298_wire_96,
Circuit298_wire_97,
Circuit298_wire_98,
Circuit298_wire_99,
Circuit298_wire_100,
Circuit298_wire_101,
Circuit298_wire_102,
Circuit298_wire_103,
Circuit298_wire_104,
Circuit298_wire_105,
Circuit298_wire_106,
Circuit298_wire_107,
Circuit298_wire_108,
Circuit298_wire_109,
Circuit298_wire_110,
Circuit298_wire_111,
Circuit298_wire_112,
Circuit298_wire_113,
Circuit298_wire_114,
Circuit298_wire_115,
Circuit298_wire_116,
Circuit298_wire_117,
Circuit298_wire_118,
Circuit298_wire_119,
Circuit298_wire_120,
Circuit298_wire_121,
Circuit298_wire_122,
Circuit298_wire_123,
Circuit298_wire_124,
Circuit298_wire_125,
Circuit298_wire_126,
Circuit298_wire_127,
Circuit298_wire_128,
Circuit298_wire_129,
Circuit298_wire_130,
Circuit298_wire_131,
Circuit298_wire_132,
Circuit298_wire_133,
Circuit298_wire_134,
Circuit298_wire_135,
Circuit298_wire_136,
Circuit298_wire_137,
Circuit298_wire_138,
Circuit298_wire_139,
Circuit298_wire_140,
Circuit298_wire_141,
Circuit298_wire_142,
Circuit298_wire_143,
Circuit298_wire_144,
Circuit298_wire_145,
Circuit298_wire_146,
Circuit298_wire_147,
Circuit298_wire_148,
Circuit298_wire_149,
Circuit298_wire_150,
Circuit298_wire_151,
Circuit298_wire_152,
Circuit298_wire_153,
Circuit298_wire_154,
Circuit298_wire_155,
Circuit298_wire_156,
Circuit298_wire_157,
Circuit298_wire_158,
Circuit298_wire_5_0,
Circuit298_wire_5_1,
Circuit298_wire_7_0,
Circuit298_wire_7_1,
Circuit298_wire_13_0,
Circuit298_wire_13_1,
Circuit298_wire_13_2,
Circuit298_wire_21_0,
Circuit298_wire_21_1,
Circuit298_wire_23_0,
Circuit298_wire_23_1,
Circuit298_wire_26_0,
Circuit298_wire_26_1,
Circuit298_wire_26_2,
Circuit298_wire_26_3,
Circuit298_wire_26_4,
Circuit298_wire_26_5,
Circuit298_wire_26_6,
Circuit298_wire_28_0,
Circuit298_wire_28_1,
Circuit298_wire_28_2,
Circuit298_wire_28_3,
Circuit298_wire_28_4,
Circuit298_wire_28_5,
Circuit298_wire_28_6,
Circuit298_wire_28_7,
Circuit298_wire_30_0,
Circuit298_wire_30_1,
Circuit298_wire_30_2,
Circuit298_wire_30_3,
Circuit298_wire_30_4,
Circuit298_wire_30_5,
Circuit298_wire_30_6,
Circuit298_wire_30_7,
Circuit298_wire_30_8,
Circuit298_wire_32_0,
Circuit298_wire_32_1,
Circuit298_wire_32_2,
Circuit298_wire_32_3,
Circuit298_wire_32_4,
Circuit298_wire_32_5,
Circuit298_wire_34_0,
Circuit298_wire_34_1,
Circuit298_wire_34_2,
Circuit298_wire_34_3,
Circuit298_wire_34_4,
Circuit298_wire_34_5,
Circuit298_wire_34_6,
Circuit298_wire_34_7,
Circuit298_wire_34_8,
Circuit298_wire_34_9,
Circuit298_wire_34_10,
Circuit298_wire_34_11,
Circuit298_wire_36_0,
Circuit298_wire_36_1,
Circuit298_wire_36_2,
Circuit298_wire_36_3,
Circuit298_wire_36_4,
Circuit298_wire_36_5,
Circuit298_wire_36_6,
Circuit298_wire_38_0,
Circuit298_wire_38_1,
Circuit298_wire_38_2,
Circuit298_wire_38_3,
Circuit298_wire_38_4,
Circuit298_wire_38_5,
Circuit298_wire_38_6,
Circuit298_wire_38_7,
Circuit298_wire_38_8,
Circuit298_wire_40_0,
Circuit298_wire_40_1,
Circuit298_wire_40_2,
Circuit298_wire_40_3,
Circuit298_wire_40_4,
Circuit298_wire_40_5,
Circuit298_wire_40_6,
Circuit298_wire_42_0,
Circuit298_wire_42_1,
Circuit298_wire_42_2,
Circuit298_wire_42_3,
Circuit298_wire_44_0,
Circuit298_wire_44_1,
Circuit298_wire_44_2,
Circuit298_wire_44_3,
Circuit298_wire_44_4,
Circuit298_wire_44_5,
Circuit298_wire_46_0,
Circuit298_wire_46_1,
Circuit298_wire_46_2,
Circuit298_wire_50_0,
Circuit298_wire_50_1,
Circuit298_wire_50_2,
Circuit298_wire_52_0,
Circuit298_wire_52_1,
Circuit298_wire_53_0,
Circuit298_wire_53_1,
Circuit298_wire_53_2,
Circuit298_wire_53_3,
Circuit298_wire_53_4,
Circuit298_wire_53_5,
Circuit298_wire_53_6,
Circuit298_wire_53_7,
Circuit298_wire_69_0,
Circuit298_wire_69_1,
Circuit298_wire_74_0,
Circuit298_wire_74_1,
Circuit298_wire_109_0,
Circuit298_wire_109_1,
Circuit298_wire_75_0,
Circuit298_wire_75_1,
Circuit298_wire_75_2,
Circuit298_wire_75_3,
Circuit298_wire_75_4,
Circuit298_wire_132_0,
Circuit298_wire_132_1,
Circuit298_wire_132_2,
Circuit298_wire_132_3,
Circuit298_wire_132_4,
Circuit298_wire_132_5,
Circuit298_wire_132_6,
Circuit298_wire_132_7,
Circuit298_wire_157_0,
Circuit298_wire_157_1,
Circuit298_wire_152_0,
Circuit298_wire_152_1,
Clock_net_0,
g0_net_0,
g1_net_0,
g2_net_0,
g117_net_0,
g132_net_0,
g66_net_0,
g118_net_0,
g133_net_0,
g67_net_0;

pin #(4) pin_0 ({Clock, g0, g1, g2}, {Clock_net_0, g0_net_0, g1_net_0, g2_net_0});

pout #(6) pout_0 ({g117_net_0, g132_net_0, g66_net_0, g118_net_0, g133_net_0, g67_net_0}, {g117, g132, g66, g118, g133, g67});
pout #(25) pout_1 ({Circuit298_wire_2, Circuit298_wire_4, Circuit298_wire_6, Circuit298_wire_8, Circuit298_wire_10, Circuit298_wire_12, Circuit298_wire_14,
					Circuit298_wire_16, Circuit298_wire_18, Circuit298_wire_20, Circuit298_wire_22, Circuit298_wire_25, Circuit298_wire_27, Circuit298_wire_29,
					Circuit298_wire_31, Circuit298_wire_33, Circuit298_wire_35, Circuit298_wire_37, Circuit298_wire_39, Circuit298_wire_41, Circuit298_wire_43,
					Circuit298_wire_45, Circuit298_wire_47, Circuit298_wire_49, Circuit298_wire_51}, 
					{Circuit298_wire_2_out, Circuit298_wire_4_out, Circuit298_wire_6_out, Circuit298_wire_8_out, Circuit298_wire_10_out, Circuit298_wire_12_out,
					Circuit298_wire_14_out, Circuit298_wire_16_out, Circuit298_wire_18_out, Circuit298_wire_20_out, Circuit298_wire_22_out, Circuit298_wire_25_out,
					Circuit298_wire_27_out, Circuit298_wire_29_out, Circuit298_wire_31_out, Circuit298_wire_33_out, Circuit298_wire_35_out, Circuit298_wire_37_out,
					Circuit298_wire_39_out, Circuit298_wire_41_out, Circuit298_wire_43_out, Circuit298_wire_45_out, Circuit298_wire_47_out, Circuit298_wire_49_out,
					Circuit298_wire_51_out});

fanout_n #(2, 0, 0) FANOUT_1 (Circuit298_wire_5, {Circuit298_wire_5_0, Circuit298_wire_5_1});
fanout_n #(2, 0, 0) FANOUT_2 (Circuit298_wire_7, {Circuit298_wire_7_0, Circuit298_wire_7_1});
fanout_n #(3, 0, 0) FANOUT_3 (Circuit298_wire_13, {Circuit298_wire_13_0, Circuit298_wire_13_1, Circuit298_wire_13_2});
fanout_n #(2, 0, 0) FANOUT_4 (Circuit298_wire_21, {Circuit298_wire_21_0, Circuit298_wire_21_1});
fanout_n #(2, 0, 0) FANOUT_5 (Circuit298_wire_23, {Circuit298_wire_23_0, Circuit298_wire_23_1});
fanout_n #(7, 0, 0) FANOUT_6 (Circuit298_wire_26, {Circuit298_wire_26_0, Circuit298_wire_26_1, Circuit298_wire_26_2, Circuit298_wire_26_3, Circuit298_wire_26_4, Circuit298_wire_26_5, Circuit298_wire_26_6});
fanout_n #(8, 0, 0) FANOUT_7 (Circuit298_wire_28, {Circuit298_wire_28_0, Circuit298_wire_28_1, Circuit298_wire_28_2, Circuit298_wire_28_3, Circuit298_wire_28_4, Circuit298_wire_28_5, Circuit298_wire_28_6, Circuit298_wire_28_7});
fanout_n #(9, 0, 0) FANOUT_8 (Circuit298_wire_30, {Circuit298_wire_30_0, Circuit298_wire_30_1, Circuit298_wire_30_2, Circuit298_wire_30_3, Circuit298_wire_30_4, Circuit298_wire_30_5, Circuit298_wire_30_6, Circuit298_wire_30_7, Circuit298_wire_30_8});
fanout_n #(6, 0, 0) FANOUT_9 (Circuit298_wire_32, {Circuit298_wire_32_0, Circuit298_wire_32_1, Circuit298_wire_32_2, Circuit298_wire_32_3, Circuit298_wire_32_4, Circuit298_wire_32_5});
fanout_n #(12, 0, 0) FANOUT_10 (Circuit298_wire_34, {Circuit298_wire_34_0, Circuit298_wire_34_1, Circuit298_wire_34_2, Circuit298_wire_34_3, Circuit298_wire_34_4, Circuit298_wire_34_5, Circuit298_wire_34_6, Circuit298_wire_34_7, Circuit298_wire_34_8, Circuit298_wire_34_9, Circuit298_wire_34_10, Circuit298_wire_34_11});
fanout_n #(7, 0, 0) FANOUT_11 (Circuit298_wire_36, {Circuit298_wire_36_0, Circuit298_wire_36_1, Circuit298_wire_36_2, Circuit298_wire_36_3, Circuit298_wire_36_4, Circuit298_wire_36_5, Circuit298_wire_36_6});
fanout_n #(9, 0, 0) FANOUT_12 (Circuit298_wire_38, {Circuit298_wire_38_0, Circuit298_wire_38_1, Circuit298_wire_38_2, Circuit298_wire_38_3, Circuit298_wire_38_4, Circuit298_wire_38_5, Circuit298_wire_38_6, Circuit298_wire_38_7, Circuit298_wire_38_8});
fanout_n #(7, 0, 0) FANOUT_13 (Circuit298_wire_40, {Circuit298_wire_40_0, Circuit298_wire_40_1, Circuit298_wire_40_2, Circuit298_wire_40_3, Circuit298_wire_40_4, Circuit298_wire_40_5, Circuit298_wire_40_6});
fanout_n #(4, 0, 0) FANOUT_14 (Circuit298_wire_42, {Circuit298_wire_42_0, Circuit298_wire_42_1, Circuit298_wire_42_2, Circuit298_wire_42_3});
fanout_n #(6, 0, 0) FANOUT_15 (Circuit298_wire_44, {Circuit298_wire_44_0, Circuit298_wire_44_1, Circuit298_wire_44_2, Circuit298_wire_44_3, Circuit298_wire_44_4, Circuit298_wire_44_5});
fanout_n #(3, 0, 0) FANOUT_16 (Circuit298_wire_46, {Circuit298_wire_46_0, Circuit298_wire_46_1, Circuit298_wire_46_2});
fanout_n #(3, 0, 0) FANOUT_17 (Circuit298_wire_50, {Circuit298_wire_50_0, Circuit298_wire_50_1, Circuit298_wire_50_2});
fanout_n #(2, 0, 0) FANOUT_18 (Circuit298_wire_52, {Circuit298_wire_52_0, Circuit298_wire_52_1});
fanout_n #(8, 0, 0) FANOUT_19 (Circuit298_wire_53, {Circuit298_wire_53_0, Circuit298_wire_53_1, Circuit298_wire_53_2, Circuit298_wire_53_3, Circuit298_wire_53_4, Circuit298_wire_53_5, Circuit298_wire_53_6, Circuit298_wire_53_7});
fanout_n #(2, 0, 0) FANOUT_20 (Circuit298_wire_69, {Circuit298_wire_69_0, Circuit298_wire_69_1});
fanout_n #(2, 0, 0) FANOUT_21 (Circuit298_wire_74, {Circuit298_wire_74_0, Circuit298_wire_74_1});
fanout_n #(2, 0, 0) FANOUT_22 (Circuit298_wire_109, {Circuit298_wire_109_0, Circuit298_wire_109_1});
fanout_n #(5, 0, 0) FANOUT_23 (Circuit298_wire_75, {Circuit298_wire_75_0, Circuit298_wire_75_1, Circuit298_wire_75_2, Circuit298_wire_75_3, Circuit298_wire_75_4});
fanout_n #(8, 0, 0) FANOUT_24 (Circuit298_wire_132, {Circuit298_wire_132_0, Circuit298_wire_132_1, Circuit298_wire_132_2, Circuit298_wire_132_3, Circuit298_wire_132_4, Circuit298_wire_132_5, Circuit298_wire_132_6, Circuit298_wire_132_7});
fanout_n #(2, 0, 0) FANOUT_25 (Circuit298_wire_157, {Circuit298_wire_157_0, Circuit298_wire_157_1});
fanout_n #(2, 0, 0) FANOUT_26 (Circuit298_wire_152, {Circuit298_wire_152_0, Circuit298_wire_152_1});


notg #(0, 0) NOT_1 (Circuit298_wire_2, Circuit298_wire_4);
notg #(0, 0) NOT_2 (Circuit298_wire_8, Circuit298_wire_10);
notg #(0, 0) NOT_3 (Circuit298_wire_14, Circuit298_wire_16);
notg #(0, 0) NOT_4 (Circuit298_wire_18, Circuit298_wire_20);
notg #(0, 0) NOT_5 (Circuit298_wire_22, Circuit298_wire_24);
notg #(0, 0) NOT_6 (Circuit298_wire_25, Circuit298_wire_27);
notg #(0, 0) NOT_7 (Circuit298_wire_29, Circuit298_wire_31);
notg #(0, 0) NOT_8 (Circuit298_wire_33, Circuit298_wire_35);
notg #(0, 0) NOT_9 (Circuit298_wire_37, Circuit298_wire_39);
notg #(0, 0) NOT_10 (Circuit298_wire_41, Circuit298_wire_43);
notg #(0, 0) NOT_11 (Circuit298_wire_45, Circuit298_wire_47);
notg #(0, 0) NOT_12 (Circuit298_wire_49, Circuit298_wire_51);
or_n #(2, 0, 0) OR_1 (Circuit298_wire_53, {Circuit298_wire_54, Circuit298_wire_55});
and_n #(4, 0, 0) AND_1 (Circuit298_wire_56, {Circuit298_wire_53_0, Circuit298_wire_57, Circuit298_wire_58, Circuit298_wire_59});
and_n #(3, 0, 0) AND_2 (Circuit298_wire_10, {Circuit298_wire_53_1, Circuit298_wire_60, Circuit298_wire_61});
notg #(0, 0) NOT_13 (Circuit298_wire_62, Circuit298_wire_53_2);
and_n #(2, 0, 0) AND_3 (Circuit298_wire_63, {Circuit298_wire_53_3, Circuit298_wire_64});
and_n #(2, 0, 0) AND_4 (Circuit298_wire_65, {Circuit298_wire_53_4, Circuit298_wire_28_0});
notg #(0, 0) NOT_14 (Circuit298_wire_66, Circuit298_wire_53_5);
and_n #(2, 0, 0) AND_5 (Circuit298_wire_67, {Circuit298_wire_53_6, Circuit298_wire_68});
and_n #(3, 0, 0) AND_6 (Circuit298_wire_69, {Circuit298_wire_44_0, Circuit298_wire_40_0, Circuit298_wire_36_0});
and_n #(4, 0, 0) AND_7 (Circuit298_wire_70, {Circuit298_wire_44_1, Circuit298_wire_32_0, Circuit298_wire_38_0, Circuit298_wire_34_0});
and_n #(2, 0, 0) AND_8 (Circuit298_wire_71, {Circuit298_wire_44_2, Circuit298_wire_72});
and_n #(2, 0, 0) AND_9 (Circuit298_wire_73, {Circuit298_wire_44_3, Circuit298_wire_38_1});
and_n #(4, 0, 0) AND_10 (Circuit298_wire_74, {Circuit298_wire_52_0, Circuit298_wire_38_2, Circuit298_wire_34_1, Circuit298_wire_75_0});
notg #(0, 0) NOT_15 (Circuit298_wire_76, Circuit298_wire_52_1);
notg #(0, 0) NOT_16 (Circuit298_wire_77, Circuit298_wire_48);
or_n #(2, 0, 0) OR_2 (Circuit298_wire_72, {Circuit298_wire_40_1, Circuit298_wire_78});
and_n #(4, 0, 0) AND_11 (Circuit298_wire_79, {Circuit298_wire_40_2, Circuit298_wire_50_0, Circuit298_wire_34_2, Circuit298_wire_75_1});
and_n #(4, 0, 0) AND_12 (Circuit298_wire_54, {Circuit298_wire_40_3, Circuit298_wire_50_1, Circuit298_wire_34_3, Circuit298_wire_75_2});
and_n #(2, 0, 0) AND_13 (Circuit298_wire_80, {Circuit298_wire_40_4, Circuit298_wire_81});
or_n #(2, 0, 0) OR_3 (Circuit298_wire_64, {Circuit298_wire_36_1, Circuit298_wire_32_1});
and_n #(2, 0, 0) AND_14 (Circuit298_wire_82, {Circuit298_wire_36_2, Circuit298_wire_13_0});
and_n #(2, 0, 0) AND_15 (Circuit298_wire_78, {Circuit298_wire_32_2, Circuit298_wire_34_4});
and_n #(2, 0, 0) AND_16 (Circuit298_wire_83, {Circuit298_wire_32_3, Circuit298_wire_84});
notg #(0, 0) NOT_17 (Circuit298_wire_81, Circuit298_wire_28_1);
and_n #(2, 0, 0) AND_17 (Circuit298_wire_85, {Circuit298_wire_28_2, Circuit298_wire_86});
and_n #(2, 0, 0) AND_18 (Circuit298_wire_87, {Circuit298_wire_28_3, Circuit298_wire_88});
and_n #(2, 0, 0) AND_19 (Circuit298_wire_89, {Circuit298_wire_42_0, Circuit298_wire_38_3});
notg #(0, 0) NOT_18 (Circuit298_wire_90, Circuit298_wire_42_1);
and_n #(2, 0, 0) AND_20 (Circuit298_wire_91, {Circuit298_wire_42_2, Circuit298_wire_66});
notg #(0, 0) NOT_19 (Circuit298_wire_86, Circuit298_wire_15);
notg #(0, 0) NOT_20 (Circuit298_wire_92, Circuit298_wire_46_0);
and_n #(2, 0, 0) AND_21 (Circuit298_wire_93, {Circuit298_wire_46_1, Circuit298_wire_26_0});
and_n #(3, 0, 0) AND_22 (Circuit298_wire_94, {Circuit298_wire_38_4, Circuit298_wire_34_5, Circuit298_wire_30_0});
notg #(0, 0) NOT_21 (Circuit298_wire_95, Circuit298_wire_34_6);
and_n #(2, 0, 0) AND_23 (Circuit298_wire_96, {Circuit298_wire_34_7, Circuit298_wire_97});
notg #(0, 0) NOT_22 (Circuit298_wire_98, Circuit298_wire_34_8);
and_n #(2, 0, 0) AND_24 (Circuit298_wire_99, {Circuit298_wire_34_9, Circuit298_wire_30_1});
and_n #(2, 0, 0) AND_25 (Circuit298_wire_100, {Circuit298_wire_30_2, Circuit298_wire_101});
notg #(0, 0) NOT_23 (Circuit298_wire_97, Circuit298_wire_30_3);
or_n #(2, 0, 0) OR_4 (Circuit298_wire_57, {Circuit298_wire_30_4, Circuit298_wire_5_0});
notg #(0, 0) NOT_24 (Circuit298_wire_102, Circuit298_wire_30_5);
notg #(0, 0) NOT_25 (Circuit298_wire_103, Circuit298_wire_30_6);
notg #(0, 0) NOT_26 (Circuit298_wire_104, Circuit298_wire_26_1);
or_n #(2, 0, 0) OR_5 (Circuit298_wire_84, {Circuit298_wire_26_2, Circuit298_wire_19});
or_n #(2, 0, 0) OR_6 (Circuit298_wire_105, {Circuit298_wire_26_3, Circuit298_wire_13_1});
and_n #(2, 0, 0) AND_26 (Circuit298_wire_106, {Circuit298_wire_23_0, Circuit298_wire_107});
and_n #(2, 0, 0) AND_27 (Circuit298_wire_55, {Circuit298_wire_23_1, Circuit298_wire_108});
nor_n #(4, 0, 0) NOR_1 (Circuit298_wire_109, {Circuit298_wire_36_3, Circuit298_wire_32_4, Circuit298_wire_26_4, Circuit298_wire_40_5});
notg #(0, 0) NOT_27 (Circuit298_wire_58, Circuit298_wire_109_0);
or_n #(2, 0, 0) OR_7 (Circuit298_wire_110, {Circuit298_wire_109_1, Circuit298_wire_83});
nor_n #(2, 0, 0) NOR_2 (Circuit298_wire_75, {Circuit298_wire_28_4, Circuit298_wire_30_7});
notg #(0, 0) NOT_28 (Circuit298_wire_59, Circuit298_wire_75_3);
notg #(0, 0) NOT_29 (Circuit298_wire_111, Circuit298_wire_75_4);
and_n #(2, 0, 0) AND_28 (Circuit298_wire_4, {Circuit298_wire_56, Circuit298_wire_112});
nand_n #(3, 0, 0) NAND_1 (Circuit298_wire_112, {Circuit298_wire_28_5, Circuit298_wire_36_4, Circuit298_wire_3});
nor_n #(3, 0, 0) NOR_3 (Circuit298_wire_113, {Circuit298_wire_32_5, Circuit298_wire_36_5, Circuit298_wire_38_5});
notg #(0, 0) NOT_30 (Circuit298_wire_114, Circuit298_wire_113);
or_n #(2, 0, 0) OR_8 (Circuit298_wire_6, {Circuit298_wire_115, Circuit298_wire_116});
and_n #(2, 0, 0) AND_29 (Circuit298_wire_116, {Circuit298_wire_65, Circuit298_wire_117});
or_n #(2, 0, 0) OR_9 (Circuit298_wire_118, {Circuit298_wire_99, Circuit298_wire_7_0});
and_n #(2, 0, 0) AND_30 (Circuit298_wire_117, {Circuit298_wire_114, Circuit298_wire_118});
nor_n #(2, 0, 0) NOR_4 (Circuit298_wire_115, {Circuit298_wire_53_7, Circuit298_wire_44_4});
nor_n #(2, 0, 0) NOR_5 (Circuit298_wire_119, {Circuit298_wire_34_10, Circuit298_wire_26_5});
or_n #(2, 0, 0) OR_10 (Circuit298_wire_61, {Circuit298_wire_102, Circuit298_wire_119});
nand_n #(2, 0, 0) NAND_2 (Circuit298_wire_60, {Circuit298_wire_28_6, Circuit298_wire_9});
or_n #(2, 0, 0) OR_11 (Circuit298_wire_12, {Circuit298_wire_67, Circuit298_wire_91});
or_n #(2, 0, 0) OR_12 (Circuit298_wire_88, {Circuit298_wire_82, Circuit298_wire_94});
or_n #(2, 0, 0) OR_13 (Circuit298_wire_68, {Circuit298_wire_120, Circuit298_wire_87});
and_n #(2, 0, 0) AND_31 (Circuit298_wire_120, {Circuit298_wire_105, Circuit298_wire_103});
and_n #(2, 0, 0) AND_32 (Circuit298_wire_16, {Circuit298_wire_63, Circuit298_wire_121});
and_n #(2, 0, 0) AND_33 (Circuit298_wire_121, {Circuit298_wire_111, Circuit298_wire_122});
or_n #(2, 0, 0) OR_14 (Circuit298_wire_122, {Circuit298_wire_80, Circuit298_wire_85});
notg #(0, 0) NOT_31 (Circuit298_wire_20, Circuit298_wire_123);
or_n #(2, 0, 0) OR_15 (Circuit298_wire_123, {Circuit298_wire_110, Circuit298_wire_124});
nor_n #(2, 0, 0) NOR_6 (Circuit298_wire_125, {Circuit298_wire_26_6, Circuit298_wire_21_0});
or_n #(2, 0, 0) OR_16 (Circuit298_wire_126, {Circuit298_wire_125, Circuit298_wire_127});
and_n #(2, 0, 0) AND_34 (Circuit298_wire_128, {Circuit298_wire_126, Circuit298_wire_98});
or_n #(2, 0, 0) OR_17 (Circuit298_wire_124, {Circuit298_wire_128, Circuit298_wire_62});
nor_n #(2, 0, 0) NOR_7 (Circuit298_wire_127, {Circuit298_wire_28_7, Circuit298_wire_38_6});
notg #(0, 0) NOT_32 (Circuit298_wire_108, Circuit298_wire_74_0);
notg #(0, 0) NOT_33 (Circuit298_wire_27, Circuit298_wire_129);
or_n #(3, 0, 0) OR_18 (Circuit298_wire_129, {Circuit298_wire_130, Circuit298_wire_131, Circuit298_wire_132_0});
and_n #(2, 0, 0) AND_35 (Circuit298_wire_133, {Circuit298_wire_73, Circuit298_wire_96});
or_n #(2, 0, 0) OR_19 (Circuit298_wire_134, {Circuit298_wire_92, Circuit298_wire_133});
and_n #(2, 0, 0) AND_36 (Circuit298_wire_130, {Circuit298_wire_134, Circuit298_wire_104});
and_n #(2, 0, 0) AND_37 (Circuit298_wire_131, {Circuit298_wire_93, Circuit298_wire_135});
notg #(0, 0) NOT_34 (Circuit298_wire_135, Circuit298_wire_70);
notg #(0, 0) NOT_35 (Circuit298_wire_24, Circuit298_wire_136);
or_n #(3, 0, 0) OR_20 (Circuit298_wire_136, {Circuit298_wire_79, Circuit298_wire_106, Circuit298_wire_132_1});
notg #(0, 0) NOT_36 (Circuit298_wire_107, Circuit298_wire_74_1);
nor_n #(2, 0, 0) NOR_8 (Circuit298_wire_43, {Circuit298_wire_44_5, Circuit298_wire_132_2});
notg #(0, 0) NOT_37 (Circuit298_wire_39, Circuit298_wire_137);
or_n #(2, 0, 0) OR_21 (Circuit298_wire_137, {Circuit298_wire_138, Circuit298_wire_71});
or_n #(2, 0, 0) OR_22 (Circuit298_wire_138, {Circuit298_wire_89, Circuit298_wire_132_3});
and_n #(3, 0, 0) AND_38 (Circuit298_wire_35, {Circuit298_wire_139, Circuit298_wire_140, Circuit298_wire_141});
nor_n #(2, 0, 0) NOR_9 (Circuit298_wire_142, {Circuit298_wire_42_3, Circuit298_wire_38_7});
or_n #(2, 0, 0) OR_23 (Circuit298_wire_141, {Circuit298_wire_95, Circuit298_wire_142});
notg #(0, 0) NOT_38 (Circuit298_wire_139, Circuit298_wire_132_4);
notg #(0, 0) NOT_39 (Circuit298_wire_140, Circuit298_wire_69_0);
notg #(0, 0) NOT_40 (Circuit298_wire_31, Circuit298_wire_143);
or_n #(2, 0, 0) OR_24 (Circuit298_wire_143, {Circuit298_wire_144, Circuit298_wire_145});
notg #(0, 0) NOT_41 (Circuit298_wire_101, Circuit298_wire_69_1);
nor_n #(2, 0, 0) NOR_10 (Circuit298_wire_146, {Circuit298_wire_40_6, Circuit298_wire_36_6});
or_n #(2, 0, 0) OR_25 (Circuit298_wire_147, {Circuit298_wire_146, Circuit298_wire_148});
or_n #(2, 0, 0) OR_26 (Circuit298_wire_144, {Circuit298_wire_100, Circuit298_wire_132_5});
and_n #(2, 0, 0) AND_39 (Circuit298_wire_145, {Circuit298_wire_147, Circuit298_wire_90});
nor_n #(3, 0, 0) NOR_11 (Circuit298_wire_148, {Circuit298_wire_34_11, Circuit298_wire_38_8, Circuit298_wire_30_8});
and_n #(2, 0, 0) AND_40 (Circuit298_wire_51, {Circuit298_wire_149, Circuit298_wire_150});
and_n #(2, 0, 0) AND_41 (Circuit298_wire_151, {Circuit298_wire_76, Circuit298_wire_152_0});
nor_n #(2, 0, 0) NOR_12 (Circuit298_wire_153, {Circuit298_wire_50_2, Circuit298_wire_152_1});
notg #(0, 0) NOT_42 (Circuit298_wire_149, Circuit298_wire_132_6);
or_n #(2, 0, 0) OR_27 (Circuit298_wire_150, {Circuit298_wire_151, Circuit298_wire_153});
and_n #(2, 0, 0) AND_42 (Circuit298_wire_47, {Circuit298_wire_154, Circuit298_wire_155});
and_n #(2, 0, 0) AND_43 (Circuit298_wire_156, {Circuit298_wire_77, Circuit298_wire_157_0});
nor_n #(2, 0, 0) NOR_13 (Circuit298_wire_158, {Circuit298_wire_46_2, Circuit298_wire_157_1});
notg #(0, 0) NOT_43 (Circuit298_wire_154, Circuit298_wire_132_7);
or_n #(2, 0, 0) OR_28 (Circuit298_wire_155, {Circuit298_wire_156, Circuit298_wire_158});
bufg #(0, 0) BUF_1 (Circuit298_wire_1, Clock_net_0);
bufg #(0, 0) BUF_2 (Circuit298_wire_132, g0_net_0);
bufg #(0, 0) BUF_3 (Circuit298_wire_157, g1_net_0);
bufg #(0, 0) BUF_4 (g117_net_0, Circuit298_wire_13_2);
bufg #(0, 0) BUF_5 (g118_net_0, Circuit298_wire_5_1);
bufg #(0, 0) BUF_6 (g132_net_0, Circuit298_wire_17);
bufg #(0, 0) BUF_7 (g133_net_0, Circuit298_wire_7_1);
bufg #(0, 0) BUF_8 (Circuit298_wire_152, g2_net_0);
bufg #(0, 0) BUF_9 (g66_net_0, Circuit298_wire_21_1);
bufg #(0, 0) BUF_10 (g67_net_0, Circuit298_wire_11);
/*	dff DFF_1  (Circuit298_wire_3, Circuit298_wire_2, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_2  (Circuit298_wire_5, Circuit298_wire_4, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_3  (Circuit298_wire_7, Circuit298_wire_6, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_4  (Circuit298_wire_9, Circuit298_wire_8, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_5  (Circuit298_wire_11, Circuit298_wire_10, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_6  (Circuit298_wire_13, Circuit298_wire_12, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_7  (Circuit298_wire_15, Circuit298_wire_14, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_8  (Circuit298_wire_17, Circuit298_wire_16, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_9  (Circuit298_wire_19, Circuit298_wire_18, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_10 (Circuit298_wire_21, Circuit298_wire_20, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_11 (Circuit298_wire_23, Circuit298_wire_22, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_12 (Circuit298_wire_26, Circuit298_wire_25, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_13 (Circuit298_wire_28, Circuit298_wire_27, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_14 (Circuit298_wire_30, Circuit298_wire_29, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_15 (Circuit298_wire_32, Circuit298_wire_31, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_16 (Circuit298_wire_34, Circuit298_wire_33, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_17 (Circuit298_wire_36, Circuit298_wire_35, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_18 (Circuit298_wire_38, Circuit298_wire_37, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_19 (Circuit298_wire_40, Circuit298_wire_39, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_20 (Circuit298_wire_42, Circuit298_wire_41, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_21 (Circuit298_wire_44, Circuit298_wire_43, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_22 (Circuit298_wire_46, Circuit298_wire_45, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_23 (Circuit298_wire_48, Circuit298_wire_47, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_24 (Circuit298_wire_50, Circuit298_wire_49, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
	dff DFF_25 (Circuit298_wire_52, Circuit298_wire_51, Circuit298_wire_1, 1'b0, 1'b0, 1'b1, NbarT, Si, reset);
*/
endmodule
