/****************************************************************************
 *                                                                          *
 *  FLAT VERSION of HIGH-LEVEL MODEL for c7552                              *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *  Verified  by: Jonathan David Hauke (jhauke@eecs.umich.edu)              *
 *                                                                          *
 *                Oct 20, 1998                                              *
 *                                                                          *
****************************************************************************/

// Flat Verilog File 
module c7552g (
	in213, in214, in215, in216, in209, in153, in154, 
	in155, in156, in157, in158, in159, in160, in151, in219, 
	in220, in221, in222, in223, in224, in225, in226, in217, 
	in231, in232, in233, in234, in235, in236, in237, in238, 
	in135, in144, in138, in147, in66, in50, in32, in35, 
	in47, in121, in94, in97, in118, in100, in124, in127, 
	in130, in103, in23, in26, in29, in41, in1486, in1480, 
	in106, in1469, in1462, in2256, in2253, in2247, in2239, in2236, 
	in2230, in2224, in2218, in2211, in4437, in4432, in4427, in4420, 
	in4415, in4410, in4405, in4400, in4394, in3749, in3743, in3737, 
	in3729, in3723, in3717, in3711, in3705, in88, in112, in87, 
	in111, in113, in110, in109, in86, in63, in64, in85, 
	in84, in83, in65, in62, in61, in60, in79, in80, 
	in81, in59, in78, in77, in56, in55, in54, in53, 
	in73, in75, in76, in74, in166, in167, in168, in169, 
	in173, in174, in175, in176, in177, in178, in179, in180, 
	in171, in189, in190, in191, in192, in193, in194, in195, 
	in196, in187, in200, in201, in202, in203, in204, in205, 
	in206, in207, in18, in12, in9, in4526, in89, in38, 
	in4528, in211, in212, in161, in227, in239, in229, in141, 
	in115, in44, in1459, in1496, in1492, in2208, in4393, in3701, 
	in3698, in114, in2204, in1455, in82, in58, in70, in69, 
	in170, in164, in165, in181, in197, in208, in198, in199, 
	in188, in172, in162, in186, in185, in182, in183, in230, 
	in218, in152, in210, in240, in228, in184, in150, in1, 
	in163, in15, in1197, in134, in133, in5, in57, in339,
	out469, out471, out327, out330, out333, out336, out324, 
	out298, out301, out304, out307, out310, out313, out316, out319, 
	out295, out347, out350, out353, out356, out359, out362, out365, 
	out368, out344, out376, out379, out382, out385, out388, out391, 
	out394, out397, out373, out419, out422, out270, out246, out273, 
	out276, out258, out264, out249, out252, out338, out321, out370, 
	out399, out416, out414, out412, out418, out410, out408, out406, 
	out404, out440, out438, out442, out444, out446, out448, out436, 
	out480, out482, out484, out486, out488, out490, out492, out494, 
	out478, out524, out526, out528, out530, out532, out534, out536, 
	out538, out522, out544, out546, out548, out550, out552, out554, 
	out556, out558, out542, out450, out496, out540, out560, out402, 
	out289, out292, out279, out278, out2, out3, out432, out453, 
	out286, out341, out281, out284, out339);

   input
	in213, in214, in215, in216, in209, in153, in154, 
	in155, in156, in157, in158, in159, in160, in151, in219, 
	in220, in221, in222, in223, in224, in225, in226, in217, 
	in231, in232, in233, in234, in235, in236, in237, in238, 
	in135, in144, in138, in147, in66, in50, in32, in35, 
	in47, in121, in94, in97, in118, in100, in124, in127, 
	in130, in103, in23, in26, in29, in41, in1486, in1480, 
	in106, in1469, in1462, in2256, in2253, in2247, in2239, in2236, 
	in2230, in2224, in2218, in2211, in4437, in4432, in4427, in4420, 
	in4415, in4410, in4405, in4400, in4394, in3749, in3743, in3737, 
	in3729, in3723, in3717, in3711, in3705, in88, in112, in87, 
	in111, in113, in110, in109, in86, in63, in64, in85, 
	in84, in83, in65, in62, in61, in60, in79, in80, 
	in81, in59, in78, in77, in56, in55, in54, in53, 
	in73, in75, in76, in74, in166, in167, in168, in169, 
	in173, in174, in175, in176, in177, in178, in179, in180, 
	in171, in189, in190, in191, in192, in193, in194, in195, 
	in196, in187, in200, in201, in202, in203, in204, in205, 
	in206, in207, in18, in12, in9, in4526, in89, in38, 
	in4528, in211, in212, in161, in227, in239, in229, in141, 
	in115, in44, in1459, in1496, in1492, in2208, in4393, in3701, 
	in3698, in114, in2204, in1455, in82, in58, in70, in69, 
	in170, in164, in165, in181, in197, in208, in198, in199, 
	in188, in172, in162, in186, in185, in182, in183, in230, 
	in218, in152, in210, in240, in228, in184, in150, in1, 
	in163, in15, in1197, in134, in133, in5, in57, in339;

   output
	out469, out471, out327, out330, out333, out336, out324, 
	out298, out301, out304, out307, out310, out313, out316, out319, 
	out295, out347, out350, out353, out356, out359, out362, out365, 
	out368, out344, out376, out379, out382, out385, out388, out391, 
	out394, out397, out373, out419, out422, out270, out246, out273, 
	out276, out258, out264, out249, out252, out338, out321, out370, 
	out399, out416, out414, out412, out418, out410, out408, out406, 
	out404, out440, out438, out442, out444, out446, out448, out436, 
	out480, out482, out484, out486, out488, out490, out492, out494, 
	out478, out524, out526, out528, out530, out532, out534, out536, 
	out538, out522, out544, out546, out548, out550, out552, out554, 
	out556, out558, out542, out450, out496, out540, out560, out402, 
	out289, out292, out279, out278, out2, out3, out432, out453, 
	out286, out341, out281, out284, out339;

nand2 M0(in12, in9, ContBusMask);
inv M00(in18, MuxSel);
inv M1_UM1_0_MM0_Mux32_0_Mux8_0_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_0_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_0_Mux1(gnd, M1_UM1_0_MM0_Mux32_0_Mux8_0_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_0_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_0_Mux2(in41, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_0_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_0_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_0_line1, M1_UM1_0_MM0_Mux32_0_Mux8_0_line2, XAbus_0);
inv M1_UM1_0_MM0_Mux32_0_Mux8_1_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_1_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_1_Mux1(in238, M1_UM1_0_MM0_Mux32_0_Mux8_1_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_1_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_1_Mux2(in29, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_1_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_1_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_1_line1, M1_UM1_0_MM0_Mux32_0_Mux8_1_line2, XAbus_1);
inv M1_UM1_0_MM0_Mux32_0_Mux8_2_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_2_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_2_Mux1(in237, M1_UM1_0_MM0_Mux32_0_Mux8_2_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_2_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_2_Mux2(in26, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_2_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_2_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_2_line1, M1_UM1_0_MM0_Mux32_0_Mux8_2_line2, XAbus_2);
inv M1_UM1_0_MM0_Mux32_0_Mux8_3_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_3_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_3_Mux1(in236, M1_UM1_0_MM0_Mux32_0_Mux8_3_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_3_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_3_Mux2(in23, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_3_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_3_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_3_line1, M1_UM1_0_MM0_Mux32_0_Mux8_3_line2, XAbus_3);
inv M1_UM1_0_MM0_Mux32_0_Mux8_4_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_4_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_4_Mux1(in235, M1_UM1_0_MM0_Mux32_0_Mux8_4_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_4_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_4_Mux2(in103, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_4_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_4_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_4_line1, M1_UM1_0_MM0_Mux32_0_Mux8_4_line2, XAbus_4);
inv M1_UM1_0_MM0_Mux32_0_Mux8_5_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_5_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_5_Mux1(in234, M1_UM1_0_MM0_Mux32_0_Mux8_5_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_5_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_5_Mux2(in130, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_5_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_5_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_5_line1, M1_UM1_0_MM0_Mux32_0_Mux8_5_line2, XAbus_5);
inv M1_UM1_0_MM0_Mux32_0_Mux8_6_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_6_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_6_Mux1(in233, M1_UM1_0_MM0_Mux32_0_Mux8_6_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_6_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_6_Mux2(in127, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_6_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_6_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_6_line1, M1_UM1_0_MM0_Mux32_0_Mux8_6_line2, XAbus_6);
inv M1_UM1_0_MM0_Mux32_0_Mux8_7_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_7_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_7_Mux1(in232, M1_UM1_0_MM0_Mux32_0_Mux8_7_Not_ContIn, M1_UM1_0_MM0_Mux32_0_Mux8_7_line1);
and2 M1_UM1_0_MM0_Mux32_0_Mux8_7_Mux2(in124, MuxSel, M1_UM1_0_MM0_Mux32_0_Mux8_7_line2);
or2 M1_UM1_0_MM0_Mux32_0_Mux8_7_Mux3(M1_UM1_0_MM0_Mux32_0_Mux8_7_line1, M1_UM1_0_MM0_Mux32_0_Mux8_7_line2, XAbus_7);
inv M1_UM1_0_MM0_Mux32_1_Mux8_0_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_0_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_0_Mux1(in231, M1_UM1_0_MM0_Mux32_1_Mux8_0_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_0_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_0_Mux2(in100, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_0_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_0_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_0_line1, M1_UM1_0_MM0_Mux32_1_Mux8_0_line2, XAbus_8);
inv M1_UM1_0_MM0_Mux32_1_Mux8_1_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_1_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_1_Mux1(in217, M1_UM1_0_MM0_Mux32_1_Mux8_1_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_1_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_1_Mux2(in118, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_1_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_1_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_1_line1, M1_UM1_0_MM0_Mux32_1_Mux8_1_line2, XAbus_9);
inv M1_UM1_0_MM0_Mux32_1_Mux8_2_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_2_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_2_Mux1(in226, M1_UM1_0_MM0_Mux32_1_Mux8_2_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_2_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_2_Mux2(in97, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_2_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_2_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_2_line1, M1_UM1_0_MM0_Mux32_1_Mux8_2_line2, XAbus_10);
inv M1_UM1_0_MM0_Mux32_1_Mux8_3_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_3_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_3_Mux1(in225, M1_UM1_0_MM0_Mux32_1_Mux8_3_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_3_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_3_Mux2(in94, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_3_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_3_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_3_line1, M1_UM1_0_MM0_Mux32_1_Mux8_3_line2, XAbus_11);
inv M1_UM1_0_MM0_Mux32_1_Mux8_4_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_4_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_4_Mux1(in224, M1_UM1_0_MM0_Mux32_1_Mux8_4_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_4_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_4_Mux2(in121, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_4_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_4_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_4_line1, M1_UM1_0_MM0_Mux32_1_Mux8_4_line2, XAbus_12);
inv M1_UM1_0_MM0_Mux32_1_Mux8_5_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_5_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_5_Mux1(in223, M1_UM1_0_MM0_Mux32_1_Mux8_5_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_5_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_5_Mux2(in47, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_5_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_5_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_5_line1, M1_UM1_0_MM0_Mux32_1_Mux8_5_line2, XAbus_13);
inv M1_UM1_0_MM0_Mux32_1_Mux8_6_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_6_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_6_Mux1(in222, M1_UM1_0_MM0_Mux32_1_Mux8_6_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_6_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_6_Mux2(in35, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_6_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_6_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_6_line1, M1_UM1_0_MM0_Mux32_1_Mux8_6_line2, XAbus_14);
inv M1_UM1_0_MM0_Mux32_1_Mux8_7_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_7_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_7_Mux1(in221, M1_UM1_0_MM0_Mux32_1_Mux8_7_Not_ContIn, M1_UM1_0_MM0_Mux32_1_Mux8_7_line1);
and2 M1_UM1_0_MM0_Mux32_1_Mux8_7_Mux2(in32, MuxSel, M1_UM1_0_MM0_Mux32_1_Mux8_7_line2);
or2 M1_UM1_0_MM0_Mux32_1_Mux8_7_Mux3(M1_UM1_0_MM0_Mux32_1_Mux8_7_line1, M1_UM1_0_MM0_Mux32_1_Mux8_7_line2, XAbus_15);
inv M1_UM1_0_MM0_Mux32_2_Mux8_0_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_0_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_0_Mux1(in220, M1_UM1_0_MM0_Mux32_2_Mux8_0_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_0_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_0_Mux2(in50, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_0_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_0_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_0_line1, M1_UM1_0_MM0_Mux32_2_Mux8_0_line2, XAbus_16);
inv M1_UM1_0_MM0_Mux32_2_Mux8_1_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_1_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_1_Mux1(in219, M1_UM1_0_MM0_Mux32_2_Mux8_1_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_1_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_1_Mux2(in66, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_1_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_1_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_1_line1, M1_UM1_0_MM0_Mux32_2_Mux8_1_line2, XAbus_17);
inv M1_UM1_0_MM0_Mux32_2_Mux8_2_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_2_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_2_Mux1(in151, M1_UM1_0_MM0_Mux32_2_Mux8_2_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_2_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_2_Mux2(in147, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_2_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_2_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_2_line1, M1_UM1_0_MM0_Mux32_2_Mux8_2_line2, XAbus_18);
inv M1_UM1_0_MM0_Mux32_2_Mux8_3_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_3_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_3_Mux1(in160, M1_UM1_0_MM0_Mux32_2_Mux8_3_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_3_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_3_Mux2(in138, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_3_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_3_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_3_line1, M1_UM1_0_MM0_Mux32_2_Mux8_3_line2, XAbus_19);
inv M1_UM1_0_MM0_Mux32_2_Mux8_4_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_4_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_4_Mux1(in159, M1_UM1_0_MM0_Mux32_2_Mux8_4_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_4_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_4_Mux2(in144, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_4_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_4_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_4_line1, M1_UM1_0_MM0_Mux32_2_Mux8_4_line2, XAbus_20);
inv M1_UM1_0_MM0_Mux32_2_Mux8_5_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_5_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_5_Mux1(in158, M1_UM1_0_MM0_Mux32_2_Mux8_5_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_5_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_5_Mux2(in135, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_5_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_5_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_5_line1, M1_UM1_0_MM0_Mux32_2_Mux8_5_line2, XAbus_21);
inv M1_UM1_0_MM0_Mux32_2_Mux8_6_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_6_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_6_Mux1(in157, M1_UM1_0_MM0_Mux32_2_Mux8_6_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_6_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_6_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_6_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_6_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_6_line1, M1_UM1_0_MM0_Mux32_2_Mux8_6_line2, M1_UM1_0_MuxOutbus_22);
inv M1_UM1_0_MM0_Mux32_2_Mux8_7_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_7_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_7_Mux1(in156, M1_UM1_0_MM0_Mux32_2_Mux8_7_Not_ContIn, M1_UM1_0_MM0_Mux32_2_Mux8_7_line1);
and2 M1_UM1_0_MM0_Mux32_2_Mux8_7_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_2_Mux8_7_line2);
or2 M1_UM1_0_MM0_Mux32_2_Mux8_7_Mux3(M1_UM1_0_MM0_Mux32_2_Mux8_7_line1, M1_UM1_0_MM0_Mux32_2_Mux8_7_line2, M1_UM1_0_MuxOutbus_23);
inv M1_UM1_0_MM0_Mux32_3_Mux8_0_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_0_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_0_Mux1(in155, M1_UM1_0_MM0_Mux32_3_Mux8_0_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_0_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_0_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_0_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_0_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_0_line1, M1_UM1_0_MM0_Mux32_3_Mux8_0_line2, M1_UM1_0_MuxOutbus_24);
inv M1_UM1_0_MM0_Mux32_3_Mux8_1_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_1_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_1_Mux1(in154, M1_UM1_0_MM0_Mux32_3_Mux8_1_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_1_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_1_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_1_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_1_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_1_line1, M1_UM1_0_MM0_Mux32_3_Mux8_1_line2, M1_UM1_0_MuxOutbus_25);
inv M1_UM1_0_MM0_Mux32_3_Mux8_2_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_2_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_2_Mux1(in153, M1_UM1_0_MM0_Mux32_3_Mux8_2_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_2_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_2_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_2_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_2_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_2_line1, M1_UM1_0_MM0_Mux32_3_Mux8_2_line2, M1_UM1_0_MuxOutbus_26);
inv M1_UM1_0_MM0_Mux32_3_Mux8_3_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_3_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_3_Mux1(in209, M1_UM1_0_MM0_Mux32_3_Mux8_3_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_3_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_3_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_3_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_3_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_3_line1, M1_UM1_0_MM0_Mux32_3_Mux8_3_line2, M1_UM1_0_MuxOutbus_27);
inv M1_UM1_0_MM0_Mux32_3_Mux8_4_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_4_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_4_Mux1(in216, M1_UM1_0_MM0_Mux32_3_Mux8_4_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_4_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_4_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_4_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_4_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_4_line1, M1_UM1_0_MM0_Mux32_3_Mux8_4_line2, M1_UM1_0_MuxOutbus_28);
inv M1_UM1_0_MM0_Mux32_3_Mux8_5_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_5_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_5_Mux1(in215, M1_UM1_0_MM0_Mux32_3_Mux8_5_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_5_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_5_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_5_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_5_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_5_line1, M1_UM1_0_MM0_Mux32_3_Mux8_5_line2, M1_UM1_0_MuxOutbus_29);
inv M1_UM1_0_MM0_Mux32_3_Mux8_6_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_6_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_6_Mux1(in214, M1_UM1_0_MM0_Mux32_3_Mux8_6_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_6_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_6_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_6_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_6_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_6_line1, M1_UM1_0_MM0_Mux32_3_Mux8_6_line2, M1_UM1_0_MuxOutbus_30);
inv M1_UM1_0_MM0_Mux32_3_Mux8_7_Mux0(MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_7_Not_ContIn);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_7_Mux1(in213, M1_UM1_0_MM0_Mux32_3_Mux8_7_Not_ContIn, M1_UM1_0_MM0_Mux32_3_Mux8_7_line1);
and2 M1_UM1_0_MM0_Mux32_3_Mux8_7_Mux2(vdd, MuxSel, M1_UM1_0_MM0_Mux32_3_Mux8_7_line2);
or2 M1_UM1_0_MM0_Mux32_3_Mux8_7_Mux3(M1_UM1_0_MM0_Mux32_3_Mux8_7_line1, M1_UM1_0_MM0_Mux32_3_Mux8_7_line2, M1_UM1_0_MuxOutbus_31);
and2 M1_UM1_0_MM1(M1_UM1_0_MuxOutbus_22, ContBusMask, XAbus_22);
and2 M1_UM1_0_MM2(M1_UM1_0_MuxOutbus_23, ContBusMask, XAbus_23);
and2 M1_UM1_0_MM3(M1_UM1_0_MuxOutbus_24, ContBusMask, XAbus_24);
and2 M1_UM1_0_MM4(M1_UM1_0_MuxOutbus_25, ContBusMask, XAbus_25);
and2 M1_UM1_0_MM5(M1_UM1_0_MuxOutbus_26, ContBusMask, XAbus_26);
and2 M1_UM1_0_MM6(M1_UM1_0_MuxOutbus_27, ContBusMask, XAbus_27);
and2 M1_UM1_0_MM7(M1_UM1_0_MuxOutbus_28, ContBusMask, XAbus_28);
and2 M1_UM1_0_MM8(M1_UM1_0_MuxOutbus_29, ContBusMask, XAbus_29);
and2 M1_UM1_0_MM9(M1_UM1_0_MuxOutbus_30, ContBusMask, XAbus_30);
and2 M1_UM1_0_MM10(M1_UM1_0_MuxOutbus_31, ContBusMask, XAbus_31);
inv M2_UM2_0_Mux0(MuxSel, M2_UM2_0_Not_ContIn);
and2 M2_UM2_0_Mux1(gnd, M2_UM2_0_Not_ContIn, M2_UM2_0_line1);
and2 M2_UM2_0_Mux2(in3701, MuxSel, M2_UM2_0_line2);
or2 M2_UM2_0_Mux3(M2_UM2_0_line1, M2_UM2_0_line2, M2_AuxXBbus_0);
and2 M2_UM2_1(in1492, in4528, M2_AuxXBbus_32);
and2 M2_UM2_2(in1496, in4528, M2_AuxXBbus_33);
inv M2_UM2_3_Inv34_0_Inv8_0(M2_AuxXBbus_0, Not_XBbus_0);
inv M2_UM2_3_Inv34_0_Inv8_1(in3705, Not_XBbus_1);
inv M2_UM2_3_Inv34_0_Inv8_2(in3711, Not_XBbus_2);
inv M2_UM2_3_Inv34_0_Inv8_3(in3717, Not_XBbus_3);
inv M2_UM2_3_Inv34_0_Inv8_4(in3723, Not_XBbus_4);
inv M2_UM2_3_Inv34_0_Inv8_5(in3729, Not_XBbus_5);
inv M2_UM2_3_Inv34_0_Inv8_6(in3737, Not_XBbus_6);
inv M2_UM2_3_Inv34_0_Inv8_7(in3743, Not_XBbus_7);
inv M2_UM2_3_Inv34_1_Inv8_0(in3749, Not_XBbus_8);
inv M2_UM2_3_Inv34_1_Inv8_1(in4394, Not_XBbus_9);
inv M2_UM2_3_Inv34_1_Inv8_2(in4400, Not_XBbus_10);
inv M2_UM2_3_Inv34_1_Inv8_3(in4405, Not_XBbus_11);
inv M2_UM2_3_Inv34_1_Inv8_4(in4410, Not_XBbus_12);
inv M2_UM2_3_Inv34_1_Inv8_5(in4415, Not_XBbus_13);
inv M2_UM2_3_Inv34_1_Inv8_6(in4420, Not_XBbus_14);
inv M2_UM2_3_Inv34_1_Inv8_7(in4427, Not_XBbus_15);
inv M2_UM2_3_Inv34_2_Inv8_0(in4432, Not_XBbus_16);
inv M2_UM2_3_Inv34_2_Inv8_1(in4437, Not_XBbus_17);
inv M2_UM2_3_Inv34_2_Inv8_2(in2211, Not_XBbus_18);
inv M2_UM2_3_Inv34_2_Inv8_3(in2218, Not_XBbus_19);
inv M2_UM2_3_Inv34_2_Inv8_4(in2224, Not_XBbus_20);
inv M2_UM2_3_Inv34_2_Inv8_5(in2230, Not_XBbus_21);
inv M2_UM2_3_Inv34_2_Inv8_6(in2236, Not_XBbus_22);
inv M2_UM2_3_Inv34_2_Inv8_7(in2239, Not_XBbus_23);
inv M2_UM2_3_Inv34_3_Inv8_0(in2247, Not_XBbus_24);
inv M2_UM2_3_Inv34_3_Inv8_1(in2253, Not_XBbus_25);
inv M2_UM2_3_Inv34_3_Inv8_2(in2256, Not_XBbus_26);
inv M2_UM2_3_Inv34_3_Inv8_3(in1462, Not_XBbus_27);
inv M2_UM2_3_Inv34_3_Inv8_4(in1469, Not_XBbus_28);
inv M2_UM2_3_Inv34_3_Inv8_5(in106, Not_XBbus_29);
inv M2_UM2_3_Inv34_3_Inv8_6(in1480, Not_XBbus_30);
inv M2_UM2_3_Inv34_3_Inv8_7(in1486, Not_XBbus_31);
inv M2_UM2_3_Inv34_4(M2_AuxXBbus_32, Not_XBbus_32);
inv M2_UM2_3_Inv34_5(M2_AuxXBbus_33, Not_XBbus_33);
inv M3_UM3_0_Mux32_0_Mux8_0_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_0_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_0_Mux1(vdd, M3_UM3_0_Mux32_0_Mux8_0_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_0_line1);
and2 M3_UM3_0_Mux32_0_Mux8_0_Mux2(in70, MuxSel, M3_UM3_0_Mux32_0_Mux8_0_line2);
or2 M3_UM3_0_Mux32_0_Mux8_0_Mux3(M3_UM3_0_Mux32_0_Mux8_0_line1, M3_UM3_0_Mux32_0_Mux8_0_line2, YAbus_0);
inv M3_UM3_0_Mux32_0_Mux8_1_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_1_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_1_Mux1(Not_XBbus_1, M3_UM3_0_Mux32_0_Mux8_1_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_1_line1);
and2 M3_UM3_0_Mux32_0_Mux8_1_Mux2(in74, MuxSel, M3_UM3_0_Mux32_0_Mux8_1_line2);
or2 M3_UM3_0_Mux32_0_Mux8_1_Mux3(M3_UM3_0_Mux32_0_Mux8_1_line1, M3_UM3_0_Mux32_0_Mux8_1_line2, YAbus_1);
inv M3_UM3_0_Mux32_0_Mux8_2_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_2_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_2_Mux1(Not_XBbus_2, M3_UM3_0_Mux32_0_Mux8_2_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_2_line1);
and2 M3_UM3_0_Mux32_0_Mux8_2_Mux2(in76, MuxSel, M3_UM3_0_Mux32_0_Mux8_2_line2);
or2 M3_UM3_0_Mux32_0_Mux8_2_Mux3(M3_UM3_0_Mux32_0_Mux8_2_line1, M3_UM3_0_Mux32_0_Mux8_2_line2, YAbus_2);
inv M3_UM3_0_Mux32_0_Mux8_3_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_3_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_3_Mux1(Not_XBbus_3, M3_UM3_0_Mux32_0_Mux8_3_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_3_line1);
and2 M3_UM3_0_Mux32_0_Mux8_3_Mux2(in75, MuxSel, M3_UM3_0_Mux32_0_Mux8_3_line2);
or2 M3_UM3_0_Mux32_0_Mux8_3_Mux3(M3_UM3_0_Mux32_0_Mux8_3_line1, M3_UM3_0_Mux32_0_Mux8_3_line2, YAbus_3);
inv M3_UM3_0_Mux32_0_Mux8_4_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_4_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_4_Mux1(Not_XBbus_4, M3_UM3_0_Mux32_0_Mux8_4_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_4_line1);
and2 M3_UM3_0_Mux32_0_Mux8_4_Mux2(in73, MuxSel, M3_UM3_0_Mux32_0_Mux8_4_line2);
or2 M3_UM3_0_Mux32_0_Mux8_4_Mux3(M3_UM3_0_Mux32_0_Mux8_4_line1, M3_UM3_0_Mux32_0_Mux8_4_line2, YAbus_4);
inv M3_UM3_0_Mux32_0_Mux8_5_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_5_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_5_Mux1(Not_XBbus_5, M3_UM3_0_Mux32_0_Mux8_5_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_5_line1);
and2 M3_UM3_0_Mux32_0_Mux8_5_Mux2(in53, MuxSel, M3_UM3_0_Mux32_0_Mux8_5_line2);
or2 M3_UM3_0_Mux32_0_Mux8_5_Mux3(M3_UM3_0_Mux32_0_Mux8_5_line1, M3_UM3_0_Mux32_0_Mux8_5_line2, YAbus_5);
inv M3_UM3_0_Mux32_0_Mux8_6_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_6_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_6_Mux1(Not_XBbus_6, M3_UM3_0_Mux32_0_Mux8_6_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_6_line1);
and2 M3_UM3_0_Mux32_0_Mux8_6_Mux2(in54, MuxSel, M3_UM3_0_Mux32_0_Mux8_6_line2);
or2 M3_UM3_0_Mux32_0_Mux8_6_Mux3(M3_UM3_0_Mux32_0_Mux8_6_line1, M3_UM3_0_Mux32_0_Mux8_6_line2, YAbus_6);
inv M3_UM3_0_Mux32_0_Mux8_7_Mux0(MuxSel, M3_UM3_0_Mux32_0_Mux8_7_Not_ContIn);
and2 M3_UM3_0_Mux32_0_Mux8_7_Mux1(Not_XBbus_7, M3_UM3_0_Mux32_0_Mux8_7_Not_ContIn, M3_UM3_0_Mux32_0_Mux8_7_line1);
and2 M3_UM3_0_Mux32_0_Mux8_7_Mux2(in55, MuxSel, M3_UM3_0_Mux32_0_Mux8_7_line2);
or2 M3_UM3_0_Mux32_0_Mux8_7_Mux3(M3_UM3_0_Mux32_0_Mux8_7_line1, M3_UM3_0_Mux32_0_Mux8_7_line2, YAbus_7);
inv M3_UM3_0_Mux32_1_Mux8_0_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_0_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_0_Mux1(Not_XBbus_8, M3_UM3_0_Mux32_1_Mux8_0_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_0_line1);
and2 M3_UM3_0_Mux32_1_Mux8_0_Mux2(in56, MuxSel, M3_UM3_0_Mux32_1_Mux8_0_line2);
or2 M3_UM3_0_Mux32_1_Mux8_0_Mux3(M3_UM3_0_Mux32_1_Mux8_0_line1, M3_UM3_0_Mux32_1_Mux8_0_line2, YAbus_8);
inv M3_UM3_0_Mux32_1_Mux8_1_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_1_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_1_Mux1(Not_XBbus_9, M3_UM3_0_Mux32_1_Mux8_1_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_1_line1);
and2 M3_UM3_0_Mux32_1_Mux8_1_Mux2(in77, MuxSel, M3_UM3_0_Mux32_1_Mux8_1_line2);
or2 M3_UM3_0_Mux32_1_Mux8_1_Mux3(M3_UM3_0_Mux32_1_Mux8_1_line1, M3_UM3_0_Mux32_1_Mux8_1_line2, YAbus_9);
inv M3_UM3_0_Mux32_1_Mux8_2_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_2_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_2_Mux1(Not_XBbus_10, M3_UM3_0_Mux32_1_Mux8_2_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_2_line1);
and2 M3_UM3_0_Mux32_1_Mux8_2_Mux2(in78, MuxSel, M3_UM3_0_Mux32_1_Mux8_2_line2);
or2 M3_UM3_0_Mux32_1_Mux8_2_Mux3(M3_UM3_0_Mux32_1_Mux8_2_line1, M3_UM3_0_Mux32_1_Mux8_2_line2, YAbus_10);
inv M3_UM3_0_Mux32_1_Mux8_3_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_3_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_3_Mux1(Not_XBbus_11, M3_UM3_0_Mux32_1_Mux8_3_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_3_line1);
and2 M3_UM3_0_Mux32_1_Mux8_3_Mux2(in59, MuxSel, M3_UM3_0_Mux32_1_Mux8_3_line2);
or2 M3_UM3_0_Mux32_1_Mux8_3_Mux3(M3_UM3_0_Mux32_1_Mux8_3_line1, M3_UM3_0_Mux32_1_Mux8_3_line2, YAbus_11);
inv M3_UM3_0_Mux32_1_Mux8_4_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_4_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_4_Mux1(Not_XBbus_12, M3_UM3_0_Mux32_1_Mux8_4_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_4_line1);
and2 M3_UM3_0_Mux32_1_Mux8_4_Mux2(in81, MuxSel, M3_UM3_0_Mux32_1_Mux8_4_line2);
or2 M3_UM3_0_Mux32_1_Mux8_4_Mux3(M3_UM3_0_Mux32_1_Mux8_4_line1, M3_UM3_0_Mux32_1_Mux8_4_line2, YAbus_12);
inv M3_UM3_0_Mux32_1_Mux8_5_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_5_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_5_Mux1(Not_XBbus_13, M3_UM3_0_Mux32_1_Mux8_5_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_5_line1);
and2 M3_UM3_0_Mux32_1_Mux8_5_Mux2(in80, MuxSel, M3_UM3_0_Mux32_1_Mux8_5_line2);
or2 M3_UM3_0_Mux32_1_Mux8_5_Mux3(M3_UM3_0_Mux32_1_Mux8_5_line1, M3_UM3_0_Mux32_1_Mux8_5_line2, YAbus_13);
inv M3_UM3_0_Mux32_1_Mux8_6_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_6_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_6_Mux1(Not_XBbus_14, M3_UM3_0_Mux32_1_Mux8_6_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_6_line1);
and2 M3_UM3_0_Mux32_1_Mux8_6_Mux2(in79, MuxSel, M3_UM3_0_Mux32_1_Mux8_6_line2);
or2 M3_UM3_0_Mux32_1_Mux8_6_Mux3(M3_UM3_0_Mux32_1_Mux8_6_line1, M3_UM3_0_Mux32_1_Mux8_6_line2, YAbus_14);
inv M3_UM3_0_Mux32_1_Mux8_7_Mux0(MuxSel, M3_UM3_0_Mux32_1_Mux8_7_Not_ContIn);
and2 M3_UM3_0_Mux32_1_Mux8_7_Mux1(Not_XBbus_15, M3_UM3_0_Mux32_1_Mux8_7_Not_ContIn, M3_UM3_0_Mux32_1_Mux8_7_line1);
and2 M3_UM3_0_Mux32_1_Mux8_7_Mux2(in60, MuxSel, M3_UM3_0_Mux32_1_Mux8_7_line2);
or2 M3_UM3_0_Mux32_1_Mux8_7_Mux3(M3_UM3_0_Mux32_1_Mux8_7_line1, M3_UM3_0_Mux32_1_Mux8_7_line2, YAbus_15);
inv M3_UM3_0_Mux32_2_Mux8_0_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_0_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_0_Mux1(Not_XBbus_16, M3_UM3_0_Mux32_2_Mux8_0_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_0_line1);
and2 M3_UM3_0_Mux32_2_Mux8_0_Mux2(in61, MuxSel, M3_UM3_0_Mux32_2_Mux8_0_line2);
or2 M3_UM3_0_Mux32_2_Mux8_0_Mux3(M3_UM3_0_Mux32_2_Mux8_0_line1, M3_UM3_0_Mux32_2_Mux8_0_line2, YAbus_16);
inv M3_UM3_0_Mux32_2_Mux8_1_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_1_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_1_Mux1(Not_XBbus_17, M3_UM3_0_Mux32_2_Mux8_1_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_1_line1);
and2 M3_UM3_0_Mux32_2_Mux8_1_Mux2(in62, MuxSel, M3_UM3_0_Mux32_2_Mux8_1_line2);
or2 M3_UM3_0_Mux32_2_Mux8_1_Mux3(M3_UM3_0_Mux32_2_Mux8_1_line1, M3_UM3_0_Mux32_2_Mux8_1_line2, YAbus_17);
inv M3_UM3_0_Mux32_2_Mux8_2_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_2_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_2_Mux1(Not_XBbus_18, M3_UM3_0_Mux32_2_Mux8_2_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_2_line1);
and2 M3_UM3_0_Mux32_2_Mux8_2_Mux2(in65, MuxSel, M3_UM3_0_Mux32_2_Mux8_2_line2);
or2 M3_UM3_0_Mux32_2_Mux8_2_Mux3(M3_UM3_0_Mux32_2_Mux8_2_line1, M3_UM3_0_Mux32_2_Mux8_2_line2, YAbus_18);
inv M3_UM3_0_Mux32_2_Mux8_3_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_3_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_3_Mux1(Not_XBbus_19, M3_UM3_0_Mux32_2_Mux8_3_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_3_line1);
and2 M3_UM3_0_Mux32_2_Mux8_3_Mux2(in83, MuxSel, M3_UM3_0_Mux32_2_Mux8_3_line2);
or2 M3_UM3_0_Mux32_2_Mux8_3_Mux3(M3_UM3_0_Mux32_2_Mux8_3_line1, M3_UM3_0_Mux32_2_Mux8_3_line2, YAbus_19);
inv M3_UM3_0_Mux32_2_Mux8_4_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_4_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_4_Mux1(Not_XBbus_20, M3_UM3_0_Mux32_2_Mux8_4_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_4_line1);
and2 M3_UM3_0_Mux32_2_Mux8_4_Mux2(in84, MuxSel, M3_UM3_0_Mux32_2_Mux8_4_line2);
or2 M3_UM3_0_Mux32_2_Mux8_4_Mux3(M3_UM3_0_Mux32_2_Mux8_4_line1, M3_UM3_0_Mux32_2_Mux8_4_line2, YAbus_20);
inv M3_UM3_0_Mux32_2_Mux8_5_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_5_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_5_Mux1(Not_XBbus_21, M3_UM3_0_Mux32_2_Mux8_5_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_5_line1);
and2 M3_UM3_0_Mux32_2_Mux8_5_Mux2(in85, MuxSel, M3_UM3_0_Mux32_2_Mux8_5_line2);
or2 M3_UM3_0_Mux32_2_Mux8_5_Mux3(M3_UM3_0_Mux32_2_Mux8_5_line1, M3_UM3_0_Mux32_2_Mux8_5_line2, YAbus_21);
inv M3_UM3_0_Mux32_2_Mux8_6_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_6_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_6_Mux1(Not_XBbus_22, M3_UM3_0_Mux32_2_Mux8_6_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_6_line1);
and2 M3_UM3_0_Mux32_2_Mux8_6_Mux2(in64, MuxSel, M3_UM3_0_Mux32_2_Mux8_6_line2);
or2 M3_UM3_0_Mux32_2_Mux8_6_Mux3(M3_UM3_0_Mux32_2_Mux8_6_line1, M3_UM3_0_Mux32_2_Mux8_6_line2, YAbus_22);
inv M3_UM3_0_Mux32_2_Mux8_7_Mux0(MuxSel, M3_UM3_0_Mux32_2_Mux8_7_Not_ContIn);
and2 M3_UM3_0_Mux32_2_Mux8_7_Mux1(Not_XBbus_23, M3_UM3_0_Mux32_2_Mux8_7_Not_ContIn, M3_UM3_0_Mux32_2_Mux8_7_line1);
and2 M3_UM3_0_Mux32_2_Mux8_7_Mux2(in63, MuxSel, M3_UM3_0_Mux32_2_Mux8_7_line2);
or2 M3_UM3_0_Mux32_2_Mux8_7_Mux3(M3_UM3_0_Mux32_2_Mux8_7_line1, M3_UM3_0_Mux32_2_Mux8_7_line2, YAbus_23);
inv M3_UM3_0_Mux32_3_Mux8_0_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_0_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_0_Mux1(Not_XBbus_24, M3_UM3_0_Mux32_3_Mux8_0_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_0_line1);
and2 M3_UM3_0_Mux32_3_Mux8_0_Mux2(in86, MuxSel, M3_UM3_0_Mux32_3_Mux8_0_line2);
or2 M3_UM3_0_Mux32_3_Mux8_0_Mux3(M3_UM3_0_Mux32_3_Mux8_0_line1, M3_UM3_0_Mux32_3_Mux8_0_line2, YAbus_24);
inv M3_UM3_0_Mux32_3_Mux8_1_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_1_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_1_Mux1(Not_XBbus_25, M3_UM3_0_Mux32_3_Mux8_1_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_1_line1);
and2 M3_UM3_0_Mux32_3_Mux8_1_Mux2(in109, MuxSel, M3_UM3_0_Mux32_3_Mux8_1_line2);
or2 M3_UM3_0_Mux32_3_Mux8_1_Mux3(M3_UM3_0_Mux32_3_Mux8_1_line1, M3_UM3_0_Mux32_3_Mux8_1_line2, YAbus_25);
inv M3_UM3_0_Mux32_3_Mux8_2_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_2_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_2_Mux1(Not_XBbus_26, M3_UM3_0_Mux32_3_Mux8_2_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_2_line1);
and2 M3_UM3_0_Mux32_3_Mux8_2_Mux2(in110, MuxSel, M3_UM3_0_Mux32_3_Mux8_2_line2);
or2 M3_UM3_0_Mux32_3_Mux8_2_Mux3(M3_UM3_0_Mux32_3_Mux8_2_line1, M3_UM3_0_Mux32_3_Mux8_2_line2, YAbus_26);
inv M3_UM3_0_Mux32_3_Mux8_3_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_3_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_3_Mux1(Not_XBbus_27, M3_UM3_0_Mux32_3_Mux8_3_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_3_line1);
and2 M3_UM3_0_Mux32_3_Mux8_3_Mux2(in113, MuxSel, M3_UM3_0_Mux32_3_Mux8_3_line2);
or2 M3_UM3_0_Mux32_3_Mux8_3_Mux3(M3_UM3_0_Mux32_3_Mux8_3_line1, M3_UM3_0_Mux32_3_Mux8_3_line2, YAbus_27);
inv M3_UM3_0_Mux32_3_Mux8_4_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_4_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_4_Mux1(Not_XBbus_28, M3_UM3_0_Mux32_3_Mux8_4_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_4_line1);
and2 M3_UM3_0_Mux32_3_Mux8_4_Mux2(in111, MuxSel, M3_UM3_0_Mux32_3_Mux8_4_line2);
or2 M3_UM3_0_Mux32_3_Mux8_4_Mux3(M3_UM3_0_Mux32_3_Mux8_4_line1, M3_UM3_0_Mux32_3_Mux8_4_line2, YAbus_28);
inv M3_UM3_0_Mux32_3_Mux8_5_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_5_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_5_Mux1(Not_XBbus_29, M3_UM3_0_Mux32_3_Mux8_5_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_5_line1);
and2 M3_UM3_0_Mux32_3_Mux8_5_Mux2(in87, MuxSel, M3_UM3_0_Mux32_3_Mux8_5_line2);
or2 M3_UM3_0_Mux32_3_Mux8_5_Mux3(M3_UM3_0_Mux32_3_Mux8_5_line1, M3_UM3_0_Mux32_3_Mux8_5_line2, YAbus_29);
inv M3_UM3_0_Mux32_3_Mux8_6_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_6_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_6_Mux1(Not_XBbus_30, M3_UM3_0_Mux32_3_Mux8_6_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_6_line1);
and2 M3_UM3_0_Mux32_3_Mux8_6_Mux2(in112, MuxSel, M3_UM3_0_Mux32_3_Mux8_6_line2);
or2 M3_UM3_0_Mux32_3_Mux8_6_Mux3(M3_UM3_0_Mux32_3_Mux8_6_line1, M3_UM3_0_Mux32_3_Mux8_6_line2, YAbus_30);
inv M3_UM3_0_Mux32_3_Mux8_7_Mux0(MuxSel, M3_UM3_0_Mux32_3_Mux8_7_Not_ContIn);
and2 M3_UM3_0_Mux32_3_Mux8_7_Mux1(Not_XBbus_31, M3_UM3_0_Mux32_3_Mux8_7_Not_ContIn, M3_UM3_0_Mux32_3_Mux8_7_line1);
and2 M3_UM3_0_Mux32_3_Mux8_7_Mux2(in88, MuxSel, M3_UM3_0_Mux32_3_Mux8_7_line2);
or2 M3_UM3_0_Mux32_3_Mux8_7_Mux3(M3_UM3_0_Mux32_3_Mux8_7_line1, M3_UM3_0_Mux32_3_Mux8_7_line2, YAbus_31);
inv M4_UM4_0_MM0_Mux32_0_Mux8_0_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_0_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_0_Mux1(gnd, M4_UM4_0_MM0_Mux32_0_Mux8_0_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_0_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_0_Mux2(in41, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_0_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_0_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_0_line1, M4_UM4_0_MM0_Mux32_0_Mux8_0_line2, YBbus_0);
inv M4_UM4_0_MM0_Mux32_0_Mux8_1_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_1_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_1_Mux1(in207, M4_UM4_0_MM0_Mux32_0_Mux8_1_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_1_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_1_Mux2(in29, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_1_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_1_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_1_line1, M4_UM4_0_MM0_Mux32_0_Mux8_1_line2, YBbus_1);
inv M4_UM4_0_MM0_Mux32_0_Mux8_2_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_2_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_2_Mux1(in206, M4_UM4_0_MM0_Mux32_0_Mux8_2_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_2_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_2_Mux2(in26, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_2_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_2_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_2_line1, M4_UM4_0_MM0_Mux32_0_Mux8_2_line2, YBbus_2);
inv M4_UM4_0_MM0_Mux32_0_Mux8_3_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_3_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_3_Mux1(in205, M4_UM4_0_MM0_Mux32_0_Mux8_3_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_3_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_3_Mux2(in23, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_3_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_3_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_3_line1, M4_UM4_0_MM0_Mux32_0_Mux8_3_line2, YBbus_3);
inv M4_UM4_0_MM0_Mux32_0_Mux8_4_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_4_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_4_Mux1(in204, M4_UM4_0_MM0_Mux32_0_Mux8_4_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_4_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_4_Mux2(in103, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_4_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_4_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_4_line1, M4_UM4_0_MM0_Mux32_0_Mux8_4_line2, YBbus_4);
inv M4_UM4_0_MM0_Mux32_0_Mux8_5_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_5_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_5_Mux1(in203, M4_UM4_0_MM0_Mux32_0_Mux8_5_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_5_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_5_Mux2(in130, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_5_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_5_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_5_line1, M4_UM4_0_MM0_Mux32_0_Mux8_5_line2, YBbus_5);
inv M4_UM4_0_MM0_Mux32_0_Mux8_6_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_6_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_6_Mux1(in202, M4_UM4_0_MM0_Mux32_0_Mux8_6_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_6_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_6_Mux2(in127, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_6_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_6_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_6_line1, M4_UM4_0_MM0_Mux32_0_Mux8_6_line2, YBbus_6);
inv M4_UM4_0_MM0_Mux32_0_Mux8_7_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_7_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_7_Mux1(in201, M4_UM4_0_MM0_Mux32_0_Mux8_7_Not_ContIn, M4_UM4_0_MM0_Mux32_0_Mux8_7_line1);
and2 M4_UM4_0_MM0_Mux32_0_Mux8_7_Mux2(in124, MuxSel, M4_UM4_0_MM0_Mux32_0_Mux8_7_line2);
or2 M4_UM4_0_MM0_Mux32_0_Mux8_7_Mux3(M4_UM4_0_MM0_Mux32_0_Mux8_7_line1, M4_UM4_0_MM0_Mux32_0_Mux8_7_line2, YBbus_7);
inv M4_UM4_0_MM0_Mux32_1_Mux8_0_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_0_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_0_Mux1(in200, M4_UM4_0_MM0_Mux32_1_Mux8_0_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_0_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_0_Mux2(in100, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_0_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_0_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_0_line1, M4_UM4_0_MM0_Mux32_1_Mux8_0_line2, YBbus_8);
inv M4_UM4_0_MM0_Mux32_1_Mux8_1_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_1_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_1_Mux1(in187, M4_UM4_0_MM0_Mux32_1_Mux8_1_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_1_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_1_Mux2(in118, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_1_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_1_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_1_line1, M4_UM4_0_MM0_Mux32_1_Mux8_1_line2, YBbus_9);
inv M4_UM4_0_MM0_Mux32_1_Mux8_2_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_2_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_2_Mux1(in196, M4_UM4_0_MM0_Mux32_1_Mux8_2_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_2_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_2_Mux2(in97, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_2_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_2_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_2_line1, M4_UM4_0_MM0_Mux32_1_Mux8_2_line2, YBbus_10);
inv M4_UM4_0_MM0_Mux32_1_Mux8_3_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_3_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_3_Mux1(in195, M4_UM4_0_MM0_Mux32_1_Mux8_3_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_3_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_3_Mux2(in94, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_3_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_3_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_3_line1, M4_UM4_0_MM0_Mux32_1_Mux8_3_line2, YBbus_11);
inv M4_UM4_0_MM0_Mux32_1_Mux8_4_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_4_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_4_Mux1(in194, M4_UM4_0_MM0_Mux32_1_Mux8_4_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_4_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_4_Mux2(in121, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_4_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_4_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_4_line1, M4_UM4_0_MM0_Mux32_1_Mux8_4_line2, YBbus_12);
inv M4_UM4_0_MM0_Mux32_1_Mux8_5_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_5_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_5_Mux1(in193, M4_UM4_0_MM0_Mux32_1_Mux8_5_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_5_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_5_Mux2(in47, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_5_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_5_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_5_line1, M4_UM4_0_MM0_Mux32_1_Mux8_5_line2, YBbus_13);
inv M4_UM4_0_MM0_Mux32_1_Mux8_6_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_6_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_6_Mux1(in192, M4_UM4_0_MM0_Mux32_1_Mux8_6_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_6_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_6_Mux2(in35, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_6_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_6_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_6_line1, M4_UM4_0_MM0_Mux32_1_Mux8_6_line2, YBbus_14);
inv M4_UM4_0_MM0_Mux32_1_Mux8_7_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_7_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_7_Mux1(in191, M4_UM4_0_MM0_Mux32_1_Mux8_7_Not_ContIn, M4_UM4_0_MM0_Mux32_1_Mux8_7_line1);
and2 M4_UM4_0_MM0_Mux32_1_Mux8_7_Mux2(in32, MuxSel, M4_UM4_0_MM0_Mux32_1_Mux8_7_line2);
or2 M4_UM4_0_MM0_Mux32_1_Mux8_7_Mux3(M4_UM4_0_MM0_Mux32_1_Mux8_7_line1, M4_UM4_0_MM0_Mux32_1_Mux8_7_line2, YBbus_15);
inv M4_UM4_0_MM0_Mux32_2_Mux8_0_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_0_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_0_Mux1(in190, M4_UM4_0_MM0_Mux32_2_Mux8_0_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_0_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_0_Mux2(in50, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_0_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_0_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_0_line1, M4_UM4_0_MM0_Mux32_2_Mux8_0_line2, YBbus_16);
inv M4_UM4_0_MM0_Mux32_2_Mux8_1_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_1_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_1_Mux1(in189, M4_UM4_0_MM0_Mux32_2_Mux8_1_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_1_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_1_Mux2(in66, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_1_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_1_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_1_line1, M4_UM4_0_MM0_Mux32_2_Mux8_1_line2, YBbus_17);
inv M4_UM4_0_MM0_Mux32_2_Mux8_2_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_2_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_2_Mux1(in171, M4_UM4_0_MM0_Mux32_2_Mux8_2_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_2_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_2_Mux2(in147, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_2_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_2_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_2_line1, M4_UM4_0_MM0_Mux32_2_Mux8_2_line2, YBbus_18);
inv M4_UM4_0_MM0_Mux32_2_Mux8_3_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_3_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_3_Mux1(in180, M4_UM4_0_MM0_Mux32_2_Mux8_3_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_3_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_3_Mux2(in138, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_3_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_3_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_3_line1, M4_UM4_0_MM0_Mux32_2_Mux8_3_line2, YBbus_19);
inv M4_UM4_0_MM0_Mux32_2_Mux8_4_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_4_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_4_Mux1(in179, M4_UM4_0_MM0_Mux32_2_Mux8_4_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_4_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_4_Mux2(in144, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_4_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_4_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_4_line1, M4_UM4_0_MM0_Mux32_2_Mux8_4_line2, YBbus_20);
inv M4_UM4_0_MM0_Mux32_2_Mux8_5_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_5_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_5_Mux1(in178, M4_UM4_0_MM0_Mux32_2_Mux8_5_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_5_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_5_Mux2(in135, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_5_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_5_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_5_line1, M4_UM4_0_MM0_Mux32_2_Mux8_5_line2, YBbus_21);
inv M4_UM4_0_MM0_Mux32_2_Mux8_6_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_6_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_6_Mux1(in177, M4_UM4_0_MM0_Mux32_2_Mux8_6_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_6_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_6_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_6_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_6_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_6_line1, M4_UM4_0_MM0_Mux32_2_Mux8_6_line2, M4_UM4_0_MuxOutbus_22);
inv M4_UM4_0_MM0_Mux32_2_Mux8_7_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_7_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_7_Mux1(in176, M4_UM4_0_MM0_Mux32_2_Mux8_7_Not_ContIn, M4_UM4_0_MM0_Mux32_2_Mux8_7_line1);
and2 M4_UM4_0_MM0_Mux32_2_Mux8_7_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_2_Mux8_7_line2);
or2 M4_UM4_0_MM0_Mux32_2_Mux8_7_Mux3(M4_UM4_0_MM0_Mux32_2_Mux8_7_line1, M4_UM4_0_MM0_Mux32_2_Mux8_7_line2, M4_UM4_0_MuxOutbus_23);
inv M4_UM4_0_MM0_Mux32_3_Mux8_0_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_0_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_0_Mux1(in175, M4_UM4_0_MM0_Mux32_3_Mux8_0_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_0_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_0_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_0_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_0_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_0_line1, M4_UM4_0_MM0_Mux32_3_Mux8_0_line2, M4_UM4_0_MuxOutbus_24);
inv M4_UM4_0_MM0_Mux32_3_Mux8_1_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_1_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_1_Mux1(in174, M4_UM4_0_MM0_Mux32_3_Mux8_1_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_1_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_1_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_1_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_1_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_1_line1, M4_UM4_0_MM0_Mux32_3_Mux8_1_line2, M4_UM4_0_MuxOutbus_25);
inv M4_UM4_0_MM0_Mux32_3_Mux8_2_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_2_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_2_Mux1(in173, M4_UM4_0_MM0_Mux32_3_Mux8_2_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_2_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_2_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_2_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_2_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_2_line1, M4_UM4_0_MM0_Mux32_3_Mux8_2_line2, M4_UM4_0_MuxOutbus_26);
inv M4_UM4_0_MM0_Mux32_3_Mux8_3_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_3_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_3_Mux1(vdd, M4_UM4_0_MM0_Mux32_3_Mux8_3_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_3_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_3_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_3_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_3_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_3_line1, M4_UM4_0_MM0_Mux32_3_Mux8_3_line2, M4_UM4_0_MuxOutbus_27);
inv M4_UM4_0_MM0_Mux32_3_Mux8_4_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_4_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_4_Mux1(in169, M4_UM4_0_MM0_Mux32_3_Mux8_4_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_4_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_4_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_4_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_4_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_4_line1, M4_UM4_0_MM0_Mux32_3_Mux8_4_line2, M4_UM4_0_MuxOutbus_28);
inv M4_UM4_0_MM0_Mux32_3_Mux8_5_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_5_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_5_Mux1(in168, M4_UM4_0_MM0_Mux32_3_Mux8_5_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_5_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_5_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_5_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_5_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_5_line1, M4_UM4_0_MM0_Mux32_3_Mux8_5_line2, M4_UM4_0_MuxOutbus_29);
inv M4_UM4_0_MM0_Mux32_3_Mux8_6_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_6_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_6_Mux1(in167, M4_UM4_0_MM0_Mux32_3_Mux8_6_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_6_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_6_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_6_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_6_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_6_line1, M4_UM4_0_MM0_Mux32_3_Mux8_6_line2, M4_UM4_0_MuxOutbus_30);
inv M4_UM4_0_MM0_Mux32_3_Mux8_7_Mux0(MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_7_Not_ContIn);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_7_Mux1(in166, M4_UM4_0_MM0_Mux32_3_Mux8_7_Not_ContIn, M4_UM4_0_MM0_Mux32_3_Mux8_7_line1);
and2 M4_UM4_0_MM0_Mux32_3_Mux8_7_Mux2(vdd, MuxSel, M4_UM4_0_MM0_Mux32_3_Mux8_7_line2);
or2 M4_UM4_0_MM0_Mux32_3_Mux8_7_Mux3(M4_UM4_0_MM0_Mux32_3_Mux8_7_line1, M4_UM4_0_MM0_Mux32_3_Mux8_7_line2, M4_UM4_0_MuxOutbus_31);
and2 M4_UM4_0_MM1(M4_UM4_0_MuxOutbus_22, ContBusMask, YBbus_22);
and2 M4_UM4_0_MM2(M4_UM4_0_MuxOutbus_23, ContBusMask, YBbus_23);
and2 M4_UM4_0_MM3(M4_UM4_0_MuxOutbus_24, ContBusMask, YBbus_24);
and2 M4_UM4_0_MM4(M4_UM4_0_MuxOutbus_25, ContBusMask, YBbus_25);
and2 M4_UM4_0_MM5(M4_UM4_0_MuxOutbus_26, ContBusMask, YBbus_26);
and2 M4_UM4_0_MM6(M4_UM4_0_MuxOutbus_27, ContBusMask, YBbus_27);
and2 M4_UM4_0_MM7(M4_UM4_0_MuxOutbus_28, ContBusMask, YBbus_28);
and2 M4_UM4_0_MM8(M4_UM4_0_MuxOutbus_29, ContBusMask, YBbus_29);
and2 M4_UM4_0_MM9(M4_UM4_0_MuxOutbus_30, ContBusMask, YBbus_30);
and2 M4_UM4_0_MM10(M4_UM4_0_MuxOutbus_31, ContBusMask, YBbus_31);
inv M4_UM4_1(in4528, M4_NotXYBext);
or2 M4_UM4_2(M4_NotXYBext, in1455, YBbus_32);
or2 M4_UM4_3(M4_NotXYBext, in2204, YBbus_33);
and2 M5_UM5_0_GP34_0_GenProp8_0(XAbus_0, Not_XBbus_0, M5_GenXbus_0);
and2 M5_UM5_0_GP34_0_GenProp8_1(XAbus_1, Not_XBbus_1, M5_GenXbus_1);
and2 M5_UM5_0_GP34_0_GenProp8_2(XAbus_2, Not_XBbus_2, M5_GenXbus_2);
and2 M5_UM5_0_GP34_0_GenProp8_3(XAbus_3, Not_XBbus_3, M5_GenXbus_3);
and2 M5_UM5_0_GP34_0_GenProp8_4(XAbus_4, Not_XBbus_4, M5_GenXbus_4);
and2 M5_UM5_0_GP34_0_GenProp8_5(XAbus_5, Not_XBbus_5, M5_GenXbus_5);
and2 M5_UM5_0_GP34_0_GenProp8_6(XAbus_6, Not_XBbus_6, M5_GenXbus_6);
and2 M5_UM5_0_GP34_0_GenProp8_7(XAbus_7, Not_XBbus_7, M5_GenXbus_7);
inv M5_UM5_0_GP34_0_GenProp8_8_Xo0(XAbus_0, M5_UM5_0_GP34_0_GenProp8_8_NotA);
inv M5_UM5_0_GP34_0_GenProp8_8_Xo1(Not_XBbus_0, M5_UM5_0_GP34_0_GenProp8_8_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_8_Xo2(M5_UM5_0_GP34_0_GenProp8_8_NotA, Not_XBbus_0, M5_UM5_0_GP34_0_GenProp8_8_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_8_Xo3(M5_UM5_0_GP34_0_GenProp8_8_NotB, XAbus_0, M5_UM5_0_GP34_0_GenProp8_8_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_8_Xo4(M5_UM5_0_GP34_0_GenProp8_8_line2, M5_UM5_0_GP34_0_GenProp8_8_line3, PropXbus_0);
inv M5_UM5_0_GP34_0_GenProp8_9_Xo0(XAbus_1, M5_UM5_0_GP34_0_GenProp8_9_NotA);
inv M5_UM5_0_GP34_0_GenProp8_9_Xo1(Not_XBbus_1, M5_UM5_0_GP34_0_GenProp8_9_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_9_Xo2(M5_UM5_0_GP34_0_GenProp8_9_NotA, Not_XBbus_1, M5_UM5_0_GP34_0_GenProp8_9_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_9_Xo3(M5_UM5_0_GP34_0_GenProp8_9_NotB, XAbus_1, M5_UM5_0_GP34_0_GenProp8_9_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_9_Xo4(M5_UM5_0_GP34_0_GenProp8_9_line2, M5_UM5_0_GP34_0_GenProp8_9_line3, PropXbus_1);
inv M5_UM5_0_GP34_0_GenProp8_10_Xo0(XAbus_2, M5_UM5_0_GP34_0_GenProp8_10_NotA);
inv M5_UM5_0_GP34_0_GenProp8_10_Xo1(Not_XBbus_2, M5_UM5_0_GP34_0_GenProp8_10_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_10_Xo2(M5_UM5_0_GP34_0_GenProp8_10_NotA, Not_XBbus_2, M5_UM5_0_GP34_0_GenProp8_10_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_10_Xo3(M5_UM5_0_GP34_0_GenProp8_10_NotB, XAbus_2, M5_UM5_0_GP34_0_GenProp8_10_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_10_Xo4(M5_UM5_0_GP34_0_GenProp8_10_line2, M5_UM5_0_GP34_0_GenProp8_10_line3, PropXbus_2);
inv M5_UM5_0_GP34_0_GenProp8_11_Xo0(XAbus_3, M5_UM5_0_GP34_0_GenProp8_11_NotA);
inv M5_UM5_0_GP34_0_GenProp8_11_Xo1(Not_XBbus_3, M5_UM5_0_GP34_0_GenProp8_11_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_11_Xo2(M5_UM5_0_GP34_0_GenProp8_11_NotA, Not_XBbus_3, M5_UM5_0_GP34_0_GenProp8_11_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_11_Xo3(M5_UM5_0_GP34_0_GenProp8_11_NotB, XAbus_3, M5_UM5_0_GP34_0_GenProp8_11_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_11_Xo4(M5_UM5_0_GP34_0_GenProp8_11_line2, M5_UM5_0_GP34_0_GenProp8_11_line3, PropXbus_3);
inv M5_UM5_0_GP34_0_GenProp8_12_Xo0(XAbus_4, M5_UM5_0_GP34_0_GenProp8_12_NotA);
inv M5_UM5_0_GP34_0_GenProp8_12_Xo1(Not_XBbus_4, M5_UM5_0_GP34_0_GenProp8_12_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_12_Xo2(M5_UM5_0_GP34_0_GenProp8_12_NotA, Not_XBbus_4, M5_UM5_0_GP34_0_GenProp8_12_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_12_Xo3(M5_UM5_0_GP34_0_GenProp8_12_NotB, XAbus_4, M5_UM5_0_GP34_0_GenProp8_12_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_12_Xo4(M5_UM5_0_GP34_0_GenProp8_12_line2, M5_UM5_0_GP34_0_GenProp8_12_line3, PropXbus_4);
inv M5_UM5_0_GP34_0_GenProp8_13_Xo0(XAbus_5, M5_UM5_0_GP34_0_GenProp8_13_NotA);
inv M5_UM5_0_GP34_0_GenProp8_13_Xo1(Not_XBbus_5, M5_UM5_0_GP34_0_GenProp8_13_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_13_Xo2(M5_UM5_0_GP34_0_GenProp8_13_NotA, Not_XBbus_5, M5_UM5_0_GP34_0_GenProp8_13_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_13_Xo3(M5_UM5_0_GP34_0_GenProp8_13_NotB, XAbus_5, M5_UM5_0_GP34_0_GenProp8_13_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_13_Xo4(M5_UM5_0_GP34_0_GenProp8_13_line2, M5_UM5_0_GP34_0_GenProp8_13_line3, PropXbus_5);
inv M5_UM5_0_GP34_0_GenProp8_14_Xo0(XAbus_6, M5_UM5_0_GP34_0_GenProp8_14_NotA);
inv M5_UM5_0_GP34_0_GenProp8_14_Xo1(Not_XBbus_6, M5_UM5_0_GP34_0_GenProp8_14_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_14_Xo2(M5_UM5_0_GP34_0_GenProp8_14_NotA, Not_XBbus_6, M5_UM5_0_GP34_0_GenProp8_14_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_14_Xo3(M5_UM5_0_GP34_0_GenProp8_14_NotB, XAbus_6, M5_UM5_0_GP34_0_GenProp8_14_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_14_Xo4(M5_UM5_0_GP34_0_GenProp8_14_line2, M5_UM5_0_GP34_0_GenProp8_14_line3, PropXbus_6);
inv M5_UM5_0_GP34_0_GenProp8_15_Xo0(XAbus_7, M5_UM5_0_GP34_0_GenProp8_15_NotA);
inv M5_UM5_0_GP34_0_GenProp8_15_Xo1(Not_XBbus_7, M5_UM5_0_GP34_0_GenProp8_15_NotB);
nand2 M5_UM5_0_GP34_0_GenProp8_15_Xo2(M5_UM5_0_GP34_0_GenProp8_15_NotA, Not_XBbus_7, M5_UM5_0_GP34_0_GenProp8_15_line2);
nand2 M5_UM5_0_GP34_0_GenProp8_15_Xo3(M5_UM5_0_GP34_0_GenProp8_15_NotB, XAbus_7, M5_UM5_0_GP34_0_GenProp8_15_line3);
nand2 M5_UM5_0_GP34_0_GenProp8_15_Xo4(M5_UM5_0_GP34_0_GenProp8_15_line2, M5_UM5_0_GP34_0_GenProp8_15_line3, PropXbus_7);
and2 M5_UM5_0_GP34_1_GenProp8_0(XAbus_8, Not_XBbus_8, M5_GenXbus_8);
and2 M5_UM5_0_GP34_1_GenProp8_1(XAbus_9, Not_XBbus_9, M5_GenXbus_9);
and2 M5_UM5_0_GP34_1_GenProp8_2(XAbus_10, Not_XBbus_10, M5_GenXbus_10);
and2 M5_UM5_0_GP34_1_GenProp8_3(XAbus_11, Not_XBbus_11, M5_GenXbus_11);
and2 M5_UM5_0_GP34_1_GenProp8_4(XAbus_12, Not_XBbus_12, M5_GenXbus_12);
and2 M5_UM5_0_GP34_1_GenProp8_5(XAbus_13, Not_XBbus_13, M5_GenXbus_13);
and2 M5_UM5_0_GP34_1_GenProp8_6(XAbus_14, Not_XBbus_14, M5_GenXbus_14);
and2 M5_UM5_0_GP34_1_GenProp8_7(XAbus_15, Not_XBbus_15, M5_GenXbus_15);
inv M5_UM5_0_GP34_1_GenProp8_8_Xo0(XAbus_8, M5_UM5_0_GP34_1_GenProp8_8_NotA);
inv M5_UM5_0_GP34_1_GenProp8_8_Xo1(Not_XBbus_8, M5_UM5_0_GP34_1_GenProp8_8_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_8_Xo2(M5_UM5_0_GP34_1_GenProp8_8_NotA, Not_XBbus_8, M5_UM5_0_GP34_1_GenProp8_8_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_8_Xo3(M5_UM5_0_GP34_1_GenProp8_8_NotB, XAbus_8, M5_UM5_0_GP34_1_GenProp8_8_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_8_Xo4(M5_UM5_0_GP34_1_GenProp8_8_line2, M5_UM5_0_GP34_1_GenProp8_8_line3, PropXbus_8);
inv M5_UM5_0_GP34_1_GenProp8_9_Xo0(XAbus_9, M5_UM5_0_GP34_1_GenProp8_9_NotA);
inv M5_UM5_0_GP34_1_GenProp8_9_Xo1(Not_XBbus_9, M5_UM5_0_GP34_1_GenProp8_9_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_9_Xo2(M5_UM5_0_GP34_1_GenProp8_9_NotA, Not_XBbus_9, M5_UM5_0_GP34_1_GenProp8_9_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_9_Xo3(M5_UM5_0_GP34_1_GenProp8_9_NotB, XAbus_9, M5_UM5_0_GP34_1_GenProp8_9_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_9_Xo4(M5_UM5_0_GP34_1_GenProp8_9_line2, M5_UM5_0_GP34_1_GenProp8_9_line3, PropXbus_9);
inv M5_UM5_0_GP34_1_GenProp8_10_Xo0(XAbus_10, M5_UM5_0_GP34_1_GenProp8_10_NotA);
inv M5_UM5_0_GP34_1_GenProp8_10_Xo1(Not_XBbus_10, M5_UM5_0_GP34_1_GenProp8_10_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_10_Xo2(M5_UM5_0_GP34_1_GenProp8_10_NotA, Not_XBbus_10, M5_UM5_0_GP34_1_GenProp8_10_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_10_Xo3(M5_UM5_0_GP34_1_GenProp8_10_NotB, XAbus_10, M5_UM5_0_GP34_1_GenProp8_10_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_10_Xo4(M5_UM5_0_GP34_1_GenProp8_10_line2, M5_UM5_0_GP34_1_GenProp8_10_line3, PropXbus_10);
inv M5_UM5_0_GP34_1_GenProp8_11_Xo0(XAbus_11, M5_UM5_0_GP34_1_GenProp8_11_NotA);
inv M5_UM5_0_GP34_1_GenProp8_11_Xo1(Not_XBbus_11, M5_UM5_0_GP34_1_GenProp8_11_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_11_Xo2(M5_UM5_0_GP34_1_GenProp8_11_NotA, Not_XBbus_11, M5_UM5_0_GP34_1_GenProp8_11_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_11_Xo3(M5_UM5_0_GP34_1_GenProp8_11_NotB, XAbus_11, M5_UM5_0_GP34_1_GenProp8_11_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_11_Xo4(M5_UM5_0_GP34_1_GenProp8_11_line2, M5_UM5_0_GP34_1_GenProp8_11_line3, PropXbus_11);
inv M5_UM5_0_GP34_1_GenProp8_12_Xo0(XAbus_12, M5_UM5_0_GP34_1_GenProp8_12_NotA);
inv M5_UM5_0_GP34_1_GenProp8_12_Xo1(Not_XBbus_12, M5_UM5_0_GP34_1_GenProp8_12_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_12_Xo2(M5_UM5_0_GP34_1_GenProp8_12_NotA, Not_XBbus_12, M5_UM5_0_GP34_1_GenProp8_12_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_12_Xo3(M5_UM5_0_GP34_1_GenProp8_12_NotB, XAbus_12, M5_UM5_0_GP34_1_GenProp8_12_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_12_Xo4(M5_UM5_0_GP34_1_GenProp8_12_line2, M5_UM5_0_GP34_1_GenProp8_12_line3, PropXbus_12);
inv M5_UM5_0_GP34_1_GenProp8_13_Xo0(XAbus_13, M5_UM5_0_GP34_1_GenProp8_13_NotA);
inv M5_UM5_0_GP34_1_GenProp8_13_Xo1(Not_XBbus_13, M5_UM5_0_GP34_1_GenProp8_13_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_13_Xo2(M5_UM5_0_GP34_1_GenProp8_13_NotA, Not_XBbus_13, M5_UM5_0_GP34_1_GenProp8_13_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_13_Xo3(M5_UM5_0_GP34_1_GenProp8_13_NotB, XAbus_13, M5_UM5_0_GP34_1_GenProp8_13_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_13_Xo4(M5_UM5_0_GP34_1_GenProp8_13_line2, M5_UM5_0_GP34_1_GenProp8_13_line3, PropXbus_13);
inv M5_UM5_0_GP34_1_GenProp8_14_Xo0(XAbus_14, M5_UM5_0_GP34_1_GenProp8_14_NotA);
inv M5_UM5_0_GP34_1_GenProp8_14_Xo1(Not_XBbus_14, M5_UM5_0_GP34_1_GenProp8_14_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_14_Xo2(M5_UM5_0_GP34_1_GenProp8_14_NotA, Not_XBbus_14, M5_UM5_0_GP34_1_GenProp8_14_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_14_Xo3(M5_UM5_0_GP34_1_GenProp8_14_NotB, XAbus_14, M5_UM5_0_GP34_1_GenProp8_14_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_14_Xo4(M5_UM5_0_GP34_1_GenProp8_14_line2, M5_UM5_0_GP34_1_GenProp8_14_line3, PropXbus_14);
inv M5_UM5_0_GP34_1_GenProp8_15_Xo0(XAbus_15, M5_UM5_0_GP34_1_GenProp8_15_NotA);
inv M5_UM5_0_GP34_1_GenProp8_15_Xo1(Not_XBbus_15, M5_UM5_0_GP34_1_GenProp8_15_NotB);
nand2 M5_UM5_0_GP34_1_GenProp8_15_Xo2(M5_UM5_0_GP34_1_GenProp8_15_NotA, Not_XBbus_15, M5_UM5_0_GP34_1_GenProp8_15_line2);
nand2 M5_UM5_0_GP34_1_GenProp8_15_Xo3(M5_UM5_0_GP34_1_GenProp8_15_NotB, XAbus_15, M5_UM5_0_GP34_1_GenProp8_15_line3);
nand2 M5_UM5_0_GP34_1_GenProp8_15_Xo4(M5_UM5_0_GP34_1_GenProp8_15_line2, M5_UM5_0_GP34_1_GenProp8_15_line3, PropXbus_15);
and2 M5_UM5_0_GP34_2_GenProp8_0(XAbus_16, Not_XBbus_16, M5_GenXbus_16);
and2 M5_UM5_0_GP34_2_GenProp8_1(XAbus_17, Not_XBbus_17, M5_GenXbus_17);
and2 M5_UM5_0_GP34_2_GenProp8_2(XAbus_18, Not_XBbus_18, M5_GenXbus_18);
and2 M5_UM5_0_GP34_2_GenProp8_3(XAbus_19, Not_XBbus_19, M5_GenXbus_19);
and2 M5_UM5_0_GP34_2_GenProp8_4(XAbus_20, Not_XBbus_20, M5_GenXbus_20);
and2 M5_UM5_0_GP34_2_GenProp8_5(XAbus_21, Not_XBbus_21, M5_GenXbus_21);
and2 M5_UM5_0_GP34_2_GenProp8_6(XAbus_22, Not_XBbus_22, M5_GenXbus_22);
and2 M5_UM5_0_GP34_2_GenProp8_7(XAbus_23, Not_XBbus_23, M5_GenXbus_23);
inv M5_UM5_0_GP34_2_GenProp8_8_Xo0(XAbus_16, M5_UM5_0_GP34_2_GenProp8_8_NotA);
inv M5_UM5_0_GP34_2_GenProp8_8_Xo1(Not_XBbus_16, M5_UM5_0_GP34_2_GenProp8_8_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_8_Xo2(M5_UM5_0_GP34_2_GenProp8_8_NotA, Not_XBbus_16, M5_UM5_0_GP34_2_GenProp8_8_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_8_Xo3(M5_UM5_0_GP34_2_GenProp8_8_NotB, XAbus_16, M5_UM5_0_GP34_2_GenProp8_8_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_8_Xo4(M5_UM5_0_GP34_2_GenProp8_8_line2, M5_UM5_0_GP34_2_GenProp8_8_line3, PropXbus_16);
inv M5_UM5_0_GP34_2_GenProp8_9_Xo0(XAbus_17, M5_UM5_0_GP34_2_GenProp8_9_NotA);
inv M5_UM5_0_GP34_2_GenProp8_9_Xo1(Not_XBbus_17, M5_UM5_0_GP34_2_GenProp8_9_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_9_Xo2(M5_UM5_0_GP34_2_GenProp8_9_NotA, Not_XBbus_17, M5_UM5_0_GP34_2_GenProp8_9_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_9_Xo3(M5_UM5_0_GP34_2_GenProp8_9_NotB, XAbus_17, M5_UM5_0_GP34_2_GenProp8_9_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_9_Xo4(M5_UM5_0_GP34_2_GenProp8_9_line2, M5_UM5_0_GP34_2_GenProp8_9_line3, PropXbus_17);
inv M5_UM5_0_GP34_2_GenProp8_10_Xo0(XAbus_18, M5_UM5_0_GP34_2_GenProp8_10_NotA);
inv M5_UM5_0_GP34_2_GenProp8_10_Xo1(Not_XBbus_18, M5_UM5_0_GP34_2_GenProp8_10_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_10_Xo2(M5_UM5_0_GP34_2_GenProp8_10_NotA, Not_XBbus_18, M5_UM5_0_GP34_2_GenProp8_10_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_10_Xo3(M5_UM5_0_GP34_2_GenProp8_10_NotB, XAbus_18, M5_UM5_0_GP34_2_GenProp8_10_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_10_Xo4(M5_UM5_0_GP34_2_GenProp8_10_line2, M5_UM5_0_GP34_2_GenProp8_10_line3, PropXbus_18);
inv M5_UM5_0_GP34_2_GenProp8_11_Xo0(XAbus_19, M5_UM5_0_GP34_2_GenProp8_11_NotA);
inv M5_UM5_0_GP34_2_GenProp8_11_Xo1(Not_XBbus_19, M5_UM5_0_GP34_2_GenProp8_11_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_11_Xo2(M5_UM5_0_GP34_2_GenProp8_11_NotA, Not_XBbus_19, M5_UM5_0_GP34_2_GenProp8_11_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_11_Xo3(M5_UM5_0_GP34_2_GenProp8_11_NotB, XAbus_19, M5_UM5_0_GP34_2_GenProp8_11_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_11_Xo4(M5_UM5_0_GP34_2_GenProp8_11_line2, M5_UM5_0_GP34_2_GenProp8_11_line3, PropXbus_19);
inv M5_UM5_0_GP34_2_GenProp8_12_Xo0(XAbus_20, M5_UM5_0_GP34_2_GenProp8_12_NotA);
inv M5_UM5_0_GP34_2_GenProp8_12_Xo1(Not_XBbus_20, M5_UM5_0_GP34_2_GenProp8_12_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_12_Xo2(M5_UM5_0_GP34_2_GenProp8_12_NotA, Not_XBbus_20, M5_UM5_0_GP34_2_GenProp8_12_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_12_Xo3(M5_UM5_0_GP34_2_GenProp8_12_NotB, XAbus_20, M5_UM5_0_GP34_2_GenProp8_12_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_12_Xo4(M5_UM5_0_GP34_2_GenProp8_12_line2, M5_UM5_0_GP34_2_GenProp8_12_line3, PropXbus_20);
inv M5_UM5_0_GP34_2_GenProp8_13_Xo0(XAbus_21, M5_UM5_0_GP34_2_GenProp8_13_NotA);
inv M5_UM5_0_GP34_2_GenProp8_13_Xo1(Not_XBbus_21, M5_UM5_0_GP34_2_GenProp8_13_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_13_Xo2(M5_UM5_0_GP34_2_GenProp8_13_NotA, Not_XBbus_21, M5_UM5_0_GP34_2_GenProp8_13_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_13_Xo3(M5_UM5_0_GP34_2_GenProp8_13_NotB, XAbus_21, M5_UM5_0_GP34_2_GenProp8_13_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_13_Xo4(M5_UM5_0_GP34_2_GenProp8_13_line2, M5_UM5_0_GP34_2_GenProp8_13_line3, PropXbus_21);
inv M5_UM5_0_GP34_2_GenProp8_14_Xo0(XAbus_22, M5_UM5_0_GP34_2_GenProp8_14_NotA);
inv M5_UM5_0_GP34_2_GenProp8_14_Xo1(Not_XBbus_22, M5_UM5_0_GP34_2_GenProp8_14_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_14_Xo2(M5_UM5_0_GP34_2_GenProp8_14_NotA, Not_XBbus_22, M5_UM5_0_GP34_2_GenProp8_14_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_14_Xo3(M5_UM5_0_GP34_2_GenProp8_14_NotB, XAbus_22, M5_UM5_0_GP34_2_GenProp8_14_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_14_Xo4(M5_UM5_0_GP34_2_GenProp8_14_line2, M5_UM5_0_GP34_2_GenProp8_14_line3, PropXbus_22);
inv M5_UM5_0_GP34_2_GenProp8_15_Xo0(XAbus_23, M5_UM5_0_GP34_2_GenProp8_15_NotA);
inv M5_UM5_0_GP34_2_GenProp8_15_Xo1(Not_XBbus_23, M5_UM5_0_GP34_2_GenProp8_15_NotB);
nand2 M5_UM5_0_GP34_2_GenProp8_15_Xo2(M5_UM5_0_GP34_2_GenProp8_15_NotA, Not_XBbus_23, M5_UM5_0_GP34_2_GenProp8_15_line2);
nand2 M5_UM5_0_GP34_2_GenProp8_15_Xo3(M5_UM5_0_GP34_2_GenProp8_15_NotB, XAbus_23, M5_UM5_0_GP34_2_GenProp8_15_line3);
nand2 M5_UM5_0_GP34_2_GenProp8_15_Xo4(M5_UM5_0_GP34_2_GenProp8_15_line2, M5_UM5_0_GP34_2_GenProp8_15_line3, PropXbus_23);
and2 M5_UM5_0_GP34_3_GenProp8_0(XAbus_24, Not_XBbus_24, M5_GenXbus_24);
and2 M5_UM5_0_GP34_3_GenProp8_1(XAbus_25, Not_XBbus_25, M5_GenXbus_25);
and2 M5_UM5_0_GP34_3_GenProp8_2(XAbus_26, Not_XBbus_26, M5_GenXbus_26);
and2 M5_UM5_0_GP34_3_GenProp8_3(XAbus_27, Not_XBbus_27, M5_GenXbus_27);
and2 M5_UM5_0_GP34_3_GenProp8_4(XAbus_28, Not_XBbus_28, M5_GenXbus_28);
and2 M5_UM5_0_GP34_3_GenProp8_5(XAbus_29, Not_XBbus_29, M5_GenXbus_29);
and2 M5_UM5_0_GP34_3_GenProp8_6(XAbus_30, Not_XBbus_30, M5_GenXbus_30);
and2 M5_UM5_0_GP34_3_GenProp8_7(XAbus_31, Not_XBbus_31, M5_GenXbus_31);
inv M5_UM5_0_GP34_3_GenProp8_8_Xo0(XAbus_24, M5_UM5_0_GP34_3_GenProp8_8_NotA);
inv M5_UM5_0_GP34_3_GenProp8_8_Xo1(Not_XBbus_24, M5_UM5_0_GP34_3_GenProp8_8_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_8_Xo2(M5_UM5_0_GP34_3_GenProp8_8_NotA, Not_XBbus_24, M5_UM5_0_GP34_3_GenProp8_8_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_8_Xo3(M5_UM5_0_GP34_3_GenProp8_8_NotB, XAbus_24, M5_UM5_0_GP34_3_GenProp8_8_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_8_Xo4(M5_UM5_0_GP34_3_GenProp8_8_line2, M5_UM5_0_GP34_3_GenProp8_8_line3, PropXbus_24);
inv M5_UM5_0_GP34_3_GenProp8_9_Xo0(XAbus_25, M5_UM5_0_GP34_3_GenProp8_9_NotA);
inv M5_UM5_0_GP34_3_GenProp8_9_Xo1(Not_XBbus_25, M5_UM5_0_GP34_3_GenProp8_9_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_9_Xo2(M5_UM5_0_GP34_3_GenProp8_9_NotA, Not_XBbus_25, M5_UM5_0_GP34_3_GenProp8_9_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_9_Xo3(M5_UM5_0_GP34_3_GenProp8_9_NotB, XAbus_25, M5_UM5_0_GP34_3_GenProp8_9_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_9_Xo4(M5_UM5_0_GP34_3_GenProp8_9_line2, M5_UM5_0_GP34_3_GenProp8_9_line3, PropXbus_25);
inv M5_UM5_0_GP34_3_GenProp8_10_Xo0(XAbus_26, M5_UM5_0_GP34_3_GenProp8_10_NotA);
inv M5_UM5_0_GP34_3_GenProp8_10_Xo1(Not_XBbus_26, M5_UM5_0_GP34_3_GenProp8_10_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_10_Xo2(M5_UM5_0_GP34_3_GenProp8_10_NotA, Not_XBbus_26, M5_UM5_0_GP34_3_GenProp8_10_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_10_Xo3(M5_UM5_0_GP34_3_GenProp8_10_NotB, XAbus_26, M5_UM5_0_GP34_3_GenProp8_10_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_10_Xo4(M5_UM5_0_GP34_3_GenProp8_10_line2, M5_UM5_0_GP34_3_GenProp8_10_line3, PropXbus_26);
inv M5_UM5_0_GP34_3_GenProp8_11_Xo0(XAbus_27, M5_UM5_0_GP34_3_GenProp8_11_NotA);
inv M5_UM5_0_GP34_3_GenProp8_11_Xo1(Not_XBbus_27, M5_UM5_0_GP34_3_GenProp8_11_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_11_Xo2(M5_UM5_0_GP34_3_GenProp8_11_NotA, Not_XBbus_27, M5_UM5_0_GP34_3_GenProp8_11_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_11_Xo3(M5_UM5_0_GP34_3_GenProp8_11_NotB, XAbus_27, M5_UM5_0_GP34_3_GenProp8_11_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_11_Xo4(M5_UM5_0_GP34_3_GenProp8_11_line2, M5_UM5_0_GP34_3_GenProp8_11_line3, PropXbus_27);
inv M5_UM5_0_GP34_3_GenProp8_12_Xo0(XAbus_28, M5_UM5_0_GP34_3_GenProp8_12_NotA);
inv M5_UM5_0_GP34_3_GenProp8_12_Xo1(Not_XBbus_28, M5_UM5_0_GP34_3_GenProp8_12_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_12_Xo2(M5_UM5_0_GP34_3_GenProp8_12_NotA, Not_XBbus_28, M5_UM5_0_GP34_3_GenProp8_12_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_12_Xo3(M5_UM5_0_GP34_3_GenProp8_12_NotB, XAbus_28, M5_UM5_0_GP34_3_GenProp8_12_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_12_Xo4(M5_UM5_0_GP34_3_GenProp8_12_line2, M5_UM5_0_GP34_3_GenProp8_12_line3, PropXbus_28);
inv M5_UM5_0_GP34_3_GenProp8_13_Xo0(XAbus_29, M5_UM5_0_GP34_3_GenProp8_13_NotA);
inv M5_UM5_0_GP34_3_GenProp8_13_Xo1(Not_XBbus_29, M5_UM5_0_GP34_3_GenProp8_13_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_13_Xo2(M5_UM5_0_GP34_3_GenProp8_13_NotA, Not_XBbus_29, M5_UM5_0_GP34_3_GenProp8_13_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_13_Xo3(M5_UM5_0_GP34_3_GenProp8_13_NotB, XAbus_29, M5_UM5_0_GP34_3_GenProp8_13_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_13_Xo4(M5_UM5_0_GP34_3_GenProp8_13_line2, M5_UM5_0_GP34_3_GenProp8_13_line3, PropXbus_29);
inv M5_UM5_0_GP34_3_GenProp8_14_Xo0(XAbus_30, M5_UM5_0_GP34_3_GenProp8_14_NotA);
inv M5_UM5_0_GP34_3_GenProp8_14_Xo1(Not_XBbus_30, M5_UM5_0_GP34_3_GenProp8_14_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_14_Xo2(M5_UM5_0_GP34_3_GenProp8_14_NotA, Not_XBbus_30, M5_UM5_0_GP34_3_GenProp8_14_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_14_Xo3(M5_UM5_0_GP34_3_GenProp8_14_NotB, XAbus_30, M5_UM5_0_GP34_3_GenProp8_14_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_14_Xo4(M5_UM5_0_GP34_3_GenProp8_14_line2, M5_UM5_0_GP34_3_GenProp8_14_line3, PropXbus_30);
inv M5_UM5_0_GP34_3_GenProp8_15_Xo0(XAbus_31, M5_UM5_0_GP34_3_GenProp8_15_NotA);
inv M5_UM5_0_GP34_3_GenProp8_15_Xo1(Not_XBbus_31, M5_UM5_0_GP34_3_GenProp8_15_NotB);
nand2 M5_UM5_0_GP34_3_GenProp8_15_Xo2(M5_UM5_0_GP34_3_GenProp8_15_NotA, Not_XBbus_31, M5_UM5_0_GP34_3_GenProp8_15_line2);
nand2 M5_UM5_0_GP34_3_GenProp8_15_Xo3(M5_UM5_0_GP34_3_GenProp8_15_NotB, XAbus_31, M5_UM5_0_GP34_3_GenProp8_15_line3);
nand2 M5_UM5_0_GP34_3_GenProp8_15_Xo4(M5_UM5_0_GP34_3_GenProp8_15_line2, M5_UM5_0_GP34_3_GenProp8_15_line3, PropXbus_31);
and2 M5_UM5_0_GP34_4(in38, Not_XBbus_32, M5_GenXbus_32);
and2 M5_UM5_0_GP34_5(in38, Not_XBbus_33, M5_GenXbus_33);
inv M5_UM5_0_GP34_6_Xo0(in38, M5_UM5_0_GP34_6_NotA);
inv M5_UM5_0_GP34_6_Xo1(Not_XBbus_32, M5_UM5_0_GP34_6_NotB);
nand2 M5_UM5_0_GP34_6_Xo2(M5_UM5_0_GP34_6_NotA, Not_XBbus_32, M5_UM5_0_GP34_6_line2);
nand2 M5_UM5_0_GP34_6_Xo3(M5_UM5_0_GP34_6_NotB, in38, M5_UM5_0_GP34_6_line3);
nand2 M5_UM5_0_GP34_6_Xo4(M5_UM5_0_GP34_6_line2, M5_UM5_0_GP34_6_line3, PropXbus_32);
inv M5_UM5_0_GP34_7_Xo0(in38, M5_UM5_0_GP34_7_NotA);
inv M5_UM5_0_GP34_7_Xo1(Not_XBbus_33, M5_UM5_0_GP34_7_NotB);
nand2 M5_UM5_0_GP34_7_Xo2(M5_UM5_0_GP34_7_NotA, Not_XBbus_33, M5_UM5_0_GP34_7_line2);
nand2 M5_UM5_0_GP34_7_Xo3(M5_UM5_0_GP34_7_NotB, in38, M5_UM5_0_GP34_7_line3);
nand2 M5_UM5_0_GP34_7_Xo4(M5_UM5_0_GP34_7_line2, M5_UM5_0_GP34_7_line3, PropXbus_33);
or2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_0(M5_GenXbus_0, PropXbus_0, LocalCarryXCin1_0);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_Ao2_0(PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_Ao2_1(M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_line0, LocalCarryXCin0_1);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_Ao3a_0(PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_Ao3a_1(PropXbus_1, PropXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_Ao3a_2(M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line1, LocalCarryXCin1_1);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_Ao3a_0(PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_Ao3a_1(PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_Ao3a_2(M5_GenXbus_2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line1, LocalCarryXCin0_2);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_0(PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_1(PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_2(PropXbus_2, PropXbus_1, PropXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_3(M5_GenXbus_2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line2, LocalCarryXCin1_2);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_0(PropXbus_3, M5_GenXbus_2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_1(PropXbus_3, PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_2(PropXbus_3, PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_3(M5_GenXbus_3, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line2, LocalCarryXCin0_3);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_0(PropXbus_3, M5_GenXbus_2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_1(PropXbus_3, PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_2(PropXbus_3, PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_3(PropXbus_3, PropXbus_2, PropXbus_1, PropXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_4(M5_GenXbus_3, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line3, LocalCarryXCin1_3);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_0(PropXbus_4, M5_GenXbus_3, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_1(PropXbus_4, PropXbus_3, M5_GenXbus_2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line1);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_2(PropXbus_4, PropXbus_3, PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line2);
and5 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_3(PropXbus_4, PropXbus_3, PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line3);
or5 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_4(M5_GenXbus_4, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line3, LocalCarryXCin0_4);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_0(PropXbus_4, M5_GenXbus_3, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_1(PropXbus_4, PropXbus_3, M5_GenXbus_2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line1);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_2(PropXbus_4, PropXbus_3, PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line2);
and5 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_3(PropXbus_4, PropXbus_3, PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line3);
and5 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_4(PropXbus_4, PropXbus_3, PropXbus_2, PropXbus_1, PropXbus_0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line4);
or6 M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_5(M5_GenXbus_4, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line2, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line3, M5_UM5_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line4, LocalCarryXCin1_4);
or2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_0(M5_GenXbus_5, PropXbus_5, LocalCarryXCin1_5);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_1_Ao2_0(PropXbus_6, M5_GenXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_1_Ao2_1(M5_GenXbus_6, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_1_line0, LocalCarryXCin0_6);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_Ao3a_0(PropXbus_6, M5_GenXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_Ao3a_1(PropXbus_6, PropXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_Ao3a_2(M5_GenXbus_6, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line1, LocalCarryXCin1_6);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_Ao3a_0(PropXbus_7, M5_GenXbus_6, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_Ao3a_1(PropXbus_7, PropXbus_6, M5_GenXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_Ao3a_2(M5_GenXbus_7, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line1, LocalCarryXCin0_7);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_0(PropXbus_7, M5_GenXbus_6, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_1(PropXbus_7, PropXbus_6, M5_GenXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_2(PropXbus_7, PropXbus_6, PropXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_3(M5_GenXbus_7, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line2, LocalCarryXCin1_7);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_0(PropXbus_8, M5_GenXbus_7, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_1(PropXbus_8, PropXbus_7, M5_GenXbus_6, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_2(PropXbus_8, PropXbus_7, PropXbus_6, M5_GenXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_3(M5_GenXbus_8, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line2, LocalCarryXCin0_8);
and2 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_0(PropXbus_8, M5_GenXbus_7, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_1(PropXbus_8, PropXbus_7, M5_GenXbus_6, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_2(PropXbus_8, PropXbus_7, PropXbus_6, M5_GenXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_3(PropXbus_8, PropXbus_7, PropXbus_6, PropXbus_5, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_4(M5_GenXbus_8, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line3, LocalCarryXCin1_8);
or2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_0(M5_GenXbus_9, PropXbus_9, LocalCarryXCin1_9);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_Ao2_0(PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_Ao2_1(M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_line0, LocalCarryXCin0_10);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_Ao3a_0(PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_Ao3a_1(PropXbus_10, PropXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_Ao3a_2(M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line1, LocalCarryXCin1_10);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_Ao3a_0(PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_Ao3a_1(PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_Ao3a_2(M5_GenXbus_11, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line1, LocalCarryXCin0_11);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_0(PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_1(PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_2(PropXbus_11, PropXbus_10, PropXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_3(M5_GenXbus_11, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line2, LocalCarryXCin1_11);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_0(PropXbus_12, M5_GenXbus_11, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_1(PropXbus_12, PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_2(PropXbus_12, PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_3(M5_GenXbus_12, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line2, LocalCarryXCin0_12);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_0(PropXbus_12, M5_GenXbus_11, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_1(PropXbus_12, PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_2(PropXbus_12, PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_3(PropXbus_12, PropXbus_11, PropXbus_10, PropXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_4(M5_GenXbus_12, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line3, LocalCarryXCin1_12);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_0(PropXbus_13, M5_GenXbus_12, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_1(PropXbus_13, PropXbus_12, M5_GenXbus_11, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line1);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_2(PropXbus_13, PropXbus_12, PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line2);
and5 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_3(PropXbus_13, PropXbus_12, PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line3);
or5 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_4(M5_GenXbus_13, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line2, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line3, LocalCarryXCin0_13);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_0(PropXbus_13, M5_GenXbus_12, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_1(PropXbus_13, PropXbus_12, M5_GenXbus_11, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line1);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_2(PropXbus_13, PropXbus_12, PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line2);
and5 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_3(PropXbus_13, PropXbus_12, PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line3);
and5 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_4(PropXbus_13, PropXbus_12, PropXbus_11, PropXbus_10, PropXbus_9, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line4);
or6 M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_5(M5_GenXbus_13, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line2, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line3, M5_UM5_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line4, LocalCarryXCin1_13);
or2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_0(M5_GenXbus_14, PropXbus_14, LocalCarryXCin1_14);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_1_Ao2_0(PropXbus_15, M5_GenXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_1_Ao2_1(M5_GenXbus_15, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_1_line0, LocalCarryXCin0_15);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_Ao3a_0(PropXbus_15, M5_GenXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_Ao3a_1(PropXbus_15, PropXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_Ao3a_2(M5_GenXbus_15, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line1, LocalCarryXCin1_15);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_Ao3a_0(PropXbus_16, M5_GenXbus_15, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_Ao3a_1(PropXbus_16, PropXbus_15, M5_GenXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_Ao3a_2(M5_GenXbus_16, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line1, LocalCarryXCin0_16);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_0(PropXbus_16, M5_GenXbus_15, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_1(PropXbus_16, PropXbus_15, M5_GenXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_2(PropXbus_16, PropXbus_15, PropXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_3(M5_GenXbus_16, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line2, LocalCarryXCin1_16);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_0(PropXbus_17, M5_GenXbus_16, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_1(PropXbus_17, PropXbus_16, M5_GenXbus_15, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_2(PropXbus_17, PropXbus_16, PropXbus_15, M5_GenXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_3(M5_GenXbus_17, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line2, LocalCarryXCin0_17);
and2 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_0(PropXbus_17, M5_GenXbus_16, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_1(PropXbus_17, PropXbus_16, M5_GenXbus_15, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_2(PropXbus_17, PropXbus_16, PropXbus_15, M5_GenXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_3(PropXbus_17, PropXbus_16, PropXbus_15, PropXbus_14, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_4(M5_GenXbus_17, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line3, LocalCarryXCin1_17);
or2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_0(M5_GenXbus_18, PropXbus_18, LocalCarryXCin1_18);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_Ao2_0(PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_Ao2_1(M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_line0, LocalCarryXCin0_19);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_Ao3a_0(PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_Ao3a_1(PropXbus_19, PropXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_Ao3a_2(M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line1, LocalCarryXCin1_19);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_Ao3a_0(PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_Ao3a_1(PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_Ao3a_2(M5_GenXbus_20, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line1, LocalCarryXCin0_20);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_0(PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_1(PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_2(PropXbus_20, PropXbus_19, PropXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_3(M5_GenXbus_20, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line2, LocalCarryXCin1_20);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_0(PropXbus_21, M5_GenXbus_20, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_1(PropXbus_21, PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_2(PropXbus_21, PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_3(M5_GenXbus_21, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line2, LocalCarryXCin0_21);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_0(PropXbus_21, M5_GenXbus_20, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_1(PropXbus_21, PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_2(PropXbus_21, PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_3(PropXbus_21, PropXbus_20, PropXbus_19, PropXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_4(M5_GenXbus_21, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line3, LocalCarryXCin1_21);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_0(PropXbus_22, M5_GenXbus_21, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_1(PropXbus_22, PropXbus_21, M5_GenXbus_20, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line1);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_2(PropXbus_22, PropXbus_21, PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line2);
and5 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_3(PropXbus_22, PropXbus_21, PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line3);
or5 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_4(M5_GenXbus_22, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line2, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line3, LocalCarryXCin0_22);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_0(PropXbus_22, M5_GenXbus_21, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_1(PropXbus_22, PropXbus_21, M5_GenXbus_20, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line1);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_2(PropXbus_22, PropXbus_21, PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line2);
and5 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_3(PropXbus_22, PropXbus_21, PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line3);
and5 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_4(PropXbus_22, PropXbus_21, PropXbus_20, PropXbus_19, PropXbus_18, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line4);
or6 M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_5(M5_GenXbus_22, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line2, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line3, M5_UM5_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line4, LocalCarryXCin1_22);
or2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_0(M5_GenXbus_23, PropXbus_23, LocalCarryXCin1_23);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_1_Ao2_0(PropXbus_24, M5_GenXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_1_Ao2_1(M5_GenXbus_24, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_1_line0, LocalCarryXCin0_24);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_Ao3a_0(PropXbus_24, M5_GenXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_Ao3a_1(PropXbus_24, PropXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_Ao3a_2(M5_GenXbus_24, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line1, LocalCarryXCin1_24);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_Ao3a_0(PropXbus_25, M5_GenXbus_24, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_Ao3a_1(PropXbus_25, PropXbus_24, M5_GenXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_Ao3a_2(M5_GenXbus_25, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line1, LocalCarryXCin0_25);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_0(PropXbus_25, M5_GenXbus_24, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_1(PropXbus_25, PropXbus_24, M5_GenXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_2(PropXbus_25, PropXbus_24, PropXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_3(M5_GenXbus_25, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line2, LocalCarryXCin1_25);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_0(PropXbus_26, M5_GenXbus_25, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_1(PropXbus_26, PropXbus_25, M5_GenXbus_24, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_2(PropXbus_26, PropXbus_25, PropXbus_24, M5_GenXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_3(M5_GenXbus_26, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line2, LocalCarryXCin0_26);
and2 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_0(PropXbus_26, M5_GenXbus_25, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_1(PropXbus_26, PropXbus_25, M5_GenXbus_24, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_2(PropXbus_26, PropXbus_25, PropXbus_24, M5_GenXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_3(PropXbus_26, PropXbus_25, PropXbus_24, PropXbus_23, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_4(M5_GenXbus_26, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line3, LocalCarryXCin1_26);
or2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_0(M5_GenXbus_27, PropXbus_27, LocalCarryXCin1_27);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_1_Ao2_0(PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_1_line0);
or2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_1_Ao2_1(M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_1_line0, LocalCarryXCin0_28);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_Ao3a_0(PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line0);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_Ao3a_1(PropXbus_28, PropXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line1);
or3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_Ao3a_2(M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line1, LocalCarryXCin1_28);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_Ao3a_0(PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line0);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_Ao3a_1(PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line1);
or3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_Ao3a_2(M5_GenXbus_29, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line1, LocalCarryXCin0_29);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_0(PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line0);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_1(PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line1);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_2(PropXbus_29, PropXbus_28, PropXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line2);
or4 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_3(M5_GenXbus_29, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line1, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line2, LocalCarryXCin1_29);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_0(PropXbus_30, M5_GenXbus_29, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line0);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_1(PropXbus_30, PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line1);
and4 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_2(PropXbus_30, PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line2);
or4 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_3(M5_GenXbus_30, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line1, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line2, LocalCarryXCin0_30);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_0(PropXbus_30, M5_GenXbus_29, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line0);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_1(PropXbus_30, PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line1);
and4 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_2(PropXbus_30, PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line2);
and4 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_3(PropXbus_30, PropXbus_29, PropXbus_28, PropXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line3);
or5 M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_4(M5_GenXbus_30, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line1, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line2, M5_UM5_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line3, LocalCarryXCin1_30);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_1_Ao5a_0(PropXbus_31, M5_GenXbus_30, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line0);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_1_Ao5a_1(PropXbus_31, PropXbus_30, M5_GenXbus_29, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line1);
and4 M5_UM5_1_CC_0_GLC34_3_GLC5_1_Ao5a_2(PropXbus_31, PropXbus_30, PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line2);
and5 M5_UM5_1_CC_0_GLC34_3_GLC5_1_Ao5a_3(PropXbus_31, PropXbus_30, PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line3);
or5 M5_UM5_1_CC_0_GLC34_3_GLC5_1_Ao5a_4(M5_GenXbus_31, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line1, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line2, M5_UM5_1_CC_0_GLC34_3_GLC5_1_line3, LocalCarryXCin0_31);
and2 M5_UM5_1_CC_0_GLC34_3_GLC5_2_Ao6a_0(PropXbus_31, M5_GenXbus_30, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line0);
and3 M5_UM5_1_CC_0_GLC34_3_GLC5_2_Ao6a_1(PropXbus_31, PropXbus_30, M5_GenXbus_29, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line1);
and4 M5_UM5_1_CC_0_GLC34_3_GLC5_2_Ao6a_2(PropXbus_31, PropXbus_30, PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line2);
and5 M5_UM5_1_CC_0_GLC34_3_GLC5_2_Ao6a_3(PropXbus_31, PropXbus_30, PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line3);
and5 M5_UM5_1_CC_0_GLC34_3_GLC5_2_Ao6a_4(PropXbus_31, PropXbus_30, PropXbus_29, PropXbus_28, PropXbus_27, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line4);
or6 M5_UM5_1_CC_0_GLC34_3_GLC5_2_Ao6a_5(M5_GenXbus_31, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line0, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line1, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line2, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line3, M5_UM5_1_CC_0_GLC34_3_GLC5_2_line4, LocalCarryXCin1_31);
or2 M5_UM5_1_CC_0_GLC34_4_GLC2_0(M5_GenXbus_32, PropXbus_32, LocalCarryXCin1_32);
and2 M5_UM5_1_CC_0_GLC34_4_GLC2_1_Ao2_0(PropXbus_33, M5_GenXbus_32, M5_UM5_1_CC_0_GLC34_4_GLC2_1_line0);
or2 M5_UM5_1_CC_0_GLC34_4_GLC2_1_Ao2_1(M5_GenXbus_33, M5_UM5_1_CC_0_GLC34_4_GLC2_1_line0, LocalCarryXCin0_33);
and2 M5_UM5_1_CC_0_GLC34_4_GLC2_2_Ao3a_0(PropXbus_33, M5_GenXbus_32, M5_UM5_1_CC_0_GLC34_4_GLC2_2_line0);
and2 M5_UM5_1_CC_0_GLC34_4_GLC2_2_Ao3a_1(PropXbus_33, PropXbus_32, M5_UM5_1_CC_0_GLC34_4_GLC2_2_line1);
or3 M5_UM5_1_CC_0_GLC34_4_GLC2_2_Ao3a_2(M5_GenXbus_33, M5_UM5_1_CC_0_GLC34_4_GLC2_2_line0, M5_UM5_1_CC_0_GLC34_4_GLC2_2_line1, LocalCarryXCin1_33);
and5 M5_UM5_1_CC_1_CGC34_0_CBC0(PropXbus_0, PropXbus_1, PropXbus_2, PropXbus_3, PropXbus_4, M5_UM5_1_CC_1_CGC34_0_Prop4_0);
and4 M5_UM5_1_CC_1_CGC34_0_CBC1(PropXbus_5, PropXbus_6, PropXbus_7, PropXbus_8, M5_UM5_1_CC_1_CGC34_0_Prop8_5);
and5 M5_UM5_1_CC_1_CGC34_0_CBC2(PropXbus_9, PropXbus_10, PropXbus_11, PropXbus_12, PropXbus_13, M5_UM5_1_CC_1_CGC34_0_Prop13_9);
and4 M5_UM5_1_CC_1_CGC34_0_CBC3(PropXbus_14, PropXbus_15, PropXbus_16, PropXbus_17, M5_UM5_1_CC_1_CGC34_0_Prop17_14);
and5 M5_UM5_1_CC_1_CGC34_0_CBC4(PropXbus_18, PropXbus_19, PropXbus_20, PropXbus_21, PropXbus_22, M5_UM5_1_CC_1_CGC34_0_Prop22_18);
and4 M5_UM5_1_CC_1_CGC34_0_CBC5(PropXbus_23, PropXbus_24, PropXbus_25, PropXbus_26, M5_UM5_1_CC_1_CGC34_0_Prop26_23);
and5 M5_UM5_1_CC_1_CGC34_0_CBC6(PropXbus_27, PropXbus_28, PropXbus_29, PropXbus_30, PropXbus_31, M5_UM5_1_CC_1_CGC34_0_Prop31_27);
and2 M5_UM5_1_CC_1_CGC34_0_CBC7(PropXbus_32, PropXbus_33, M5_UM5_1_CC_1_CGC34_0_Prop33_32);
and2 M5_UM5_1_CC_1_CGC34_0_CBC8(M5_UM5_1_CC_1_CGC34_0_Prop4_0, M5_UM5_1_CC_1_CGC34_0_Prop8_5, M5_UM5_1_CC_1_CGC34_0_Prop8_0);
and2 M5_UM5_1_CC_1_CGC34_0_CBC9(M5_UM5_1_CC_1_CGC34_0_Prop13_9, M5_UM5_1_CC_1_CGC34_0_Prop17_14, M5_UM5_1_CC_1_CGC34_0_Prop17_9);
and2 M5_UM5_1_CC_1_CGC34_0_CBC10(M5_UM5_1_CC_1_CGC34_0_Prop22_18, M5_UM5_1_CC_1_CGC34_0_Prop26_23, M5_UM5_1_CC_1_CGC34_0_Prop26_18);
and2 M5_UM5_1_CC_1_CGC34_0_CBC11(M5_UM5_1_CC_1_CGC34_0_Prop31_27, M5_UM5_1_CC_1_CGC34_0_Prop33_32, M5_UM5_1_CC_1_CGC34_0_Prop33_27);
and2 M5_UM5_1_CC_1_CGC34_0_CBC12_Ao2_0(in4526, M5_UM5_1_CC_1_CGC34_0_Prop4_0, M5_UM5_1_CC_1_CGC34_0_CBC12_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CBC12_Ao2_1(LocalCarryXCin0_4, M5_UM5_1_CC_1_CGC34_0_CBC12_line0, CarryXbus_4);
inv M5_UM5_1_CC_1_CGC34_0_CGC13_Mux0(CarryXbus_4, M5_UM5_1_CC_1_CGC34_0_CGC13_Not_ContIn);
and2 M5_UM5_1_CC_1_CGC34_0_CGC13_Mux1(LocalCarryXCin0_8, M5_UM5_1_CC_1_CGC34_0_CGC13_Not_ContIn, M5_UM5_1_CC_1_CGC34_0_CGC13_line1);
and2 M5_UM5_1_CC_1_CGC34_0_CGC13_Mux2(LocalCarryXCin1_8, CarryXbus_4, M5_UM5_1_CC_1_CGC34_0_CGC13_line2);
or2 M5_UM5_1_CC_1_CGC34_0_CGC13_Mux3(M5_UM5_1_CC_1_CGC34_0_CGC13_line1, M5_UM5_1_CC_1_CGC34_0_CGC13_line2, CarryXbus_8);
and2 M5_UM5_1_CC_1_CGC34_0_GGC14_Ao2_0(CarryXbus_8, M5_UM5_1_CC_1_CGC34_0_Prop13_9, M5_UM5_1_CC_1_CGC34_0_GGC14_line0);
or2 M5_UM5_1_CC_1_CGC34_0_GGC14_Ao2_1(LocalCarryXCin0_13, M5_UM5_1_CC_1_CGC34_0_GGC14_line0, CarryXbus_13);
and2 M5_UM5_1_CC_1_CGC34_0_CGC15_Ao2_0(LocalCarryXCin0_13, M5_UM5_1_CC_1_CGC34_0_Prop17_14, M5_UM5_1_CC_1_CGC34_0_CGC15_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CGC15_Ao2_1(LocalCarryXCin0_17, M5_UM5_1_CC_1_CGC34_0_CGC15_line0, M5_UM5_1_CC_1_CGC34_0_LocalCarry17_9);
and2 M5_UM5_1_CC_1_CGC34_0_CGC16_Ao2_0(LocalCarryXCin0_4, M5_UM5_1_CC_1_CGC34_0_Prop8_5, M5_UM5_1_CC_1_CGC34_0_CGC16_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CGC16_Ao2_1(LocalCarryXCin0_8, M5_UM5_1_CC_1_CGC34_0_CGC16_line0, M5_UM5_1_CC_1_CGC34_0_LocalCarry8_0);
and2 M5_UM5_1_CC_1_CGC34_0_CGC17_Ao3a_0(M5_UM5_1_CC_1_CGC34_0_Prop17_9, M5_UM5_1_CC_1_CGC34_0_LocalCarry8_0, M5_UM5_1_CC_1_CGC34_0_CGC17_line0);
and3 M5_UM5_1_CC_1_CGC34_0_CGC17_Ao3a_1(M5_UM5_1_CC_1_CGC34_0_Prop17_9, M5_UM5_1_CC_1_CGC34_0_Prop8_0, in4526, M5_UM5_1_CC_1_CGC34_0_CGC17_line1);
or3 M5_UM5_1_CC_1_CGC34_0_CGC17_Ao3a_2(M5_UM5_1_CC_1_CGC34_0_LocalCarry17_9, M5_UM5_1_CC_1_CGC34_0_CGC17_line0, M5_UM5_1_CC_1_CGC34_0_CGC17_line1, CarryXbus_17);
and2 M5_UM5_1_CC_1_CGC34_0_CGC18_Ao2_0(CarryXbus_17, M5_UM5_1_CC_1_CGC34_0_Prop22_18, M5_UM5_1_CC_1_CGC34_0_CGC18_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CGC18_Ao2_1(LocalCarryXCin0_22, M5_UM5_1_CC_1_CGC34_0_CGC18_line0, CarryXbus_22);
and2 M5_UM5_1_CC_1_CGC34_0_CGC19_Ao2_0(LocalCarryXCin0_22, M5_UM5_1_CC_1_CGC34_0_Prop26_23, M5_UM5_1_CC_1_CGC34_0_CGC19_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CGC19_Ao2_1(LocalCarryXCin0_26, M5_UM5_1_CC_1_CGC34_0_CGC19_line0, M5_UM5_1_CC_1_CGC34_0_LocalCarry26_18);
and2 M5_UM5_1_CC_1_CGC34_0_CGC20_Ao4a_0(M5_UM5_1_CC_1_CGC34_0_Prop26_18, M5_UM5_1_CC_1_CGC34_0_LocalCarry17_9, M5_UM5_1_CC_1_CGC34_0_CGC20_line0);
and3 M5_UM5_1_CC_1_CGC34_0_CGC20_Ao4a_1(M5_UM5_1_CC_1_CGC34_0_Prop26_18, M5_UM5_1_CC_1_CGC34_0_Prop17_9, M5_UM5_1_CC_1_CGC34_0_LocalCarry8_0, M5_UM5_1_CC_1_CGC34_0_CGC20_line1);
and4 M5_UM5_1_CC_1_CGC34_0_CGC20_Ao4a_2(M5_UM5_1_CC_1_CGC34_0_Prop26_18, M5_UM5_1_CC_1_CGC34_0_Prop17_9, M5_UM5_1_CC_1_CGC34_0_Prop8_0, in4526, M5_UM5_1_CC_1_CGC34_0_CGC20_line2);
or4 M5_UM5_1_CC_1_CGC34_0_CGC20_Ao4a_3(M5_UM5_1_CC_1_CGC34_0_LocalCarry26_18, M5_UM5_1_CC_1_CGC34_0_CGC20_line0, M5_UM5_1_CC_1_CGC34_0_CGC20_line1, M5_UM5_1_CC_1_CGC34_0_CGC20_line2, CarryXbus_26);
and2 M5_UM5_1_CC_1_CGC34_0_CGC21_Ao2_0(CarryXbus_26, M5_UM5_1_CC_1_CGC34_0_Prop31_27, M5_UM5_1_CC_1_CGC34_0_CGC21_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CGC21_Ao2_1(LocalCarryXCin0_31, M5_UM5_1_CC_1_CGC34_0_CGC21_line0, CarryXbus_31);
and2 M5_UM5_1_CC_1_CGC34_0_CGC22_Ao2_0(LocalCarryXCin0_31, M5_UM5_1_CC_1_CGC34_0_Prop33_32, M5_UM5_1_CC_1_CGC34_0_CGC22_line0);
or2 M5_UM5_1_CC_1_CGC34_0_CGC22_Ao2_1(LocalCarryXCin0_33, M5_UM5_1_CC_1_CGC34_0_CGC22_line0, M5_UM5_1_CC_1_CGC34_0_LocalCarry33_27);
and2 M5_UM5_1_CC_1_CGC34_0_CGC23_Ao5a_0(M5_UM5_1_CC_1_CGC34_0_Prop33_27, M5_UM5_1_CC_1_CGC34_0_LocalCarry26_18, M5_UM5_1_CC_1_CGC34_0_CGC23_line0);
and3 M5_UM5_1_CC_1_CGC34_0_CGC23_Ao5a_1(M5_UM5_1_CC_1_CGC34_0_Prop33_27, M5_UM5_1_CC_1_CGC34_0_Prop26_18, M5_UM5_1_CC_1_CGC34_0_LocalCarry17_9, M5_UM5_1_CC_1_CGC34_0_CGC23_line1);
and4 M5_UM5_1_CC_1_CGC34_0_CGC23_Ao5a_2(M5_UM5_1_CC_1_CGC34_0_Prop33_27, M5_UM5_1_CC_1_CGC34_0_Prop26_18, M5_UM5_1_CC_1_CGC34_0_Prop17_9, M5_UM5_1_CC_1_CGC34_0_LocalCarry8_0, M5_UM5_1_CC_1_CGC34_0_CGC23_line2);
and5 M5_UM5_1_CC_1_CGC34_0_CGC23_Ao5a_3(M5_UM5_1_CC_1_CGC34_0_Prop33_27, M5_UM5_1_CC_1_CGC34_0_Prop26_18, M5_UM5_1_CC_1_CGC34_0_Prop17_9, M5_UM5_1_CC_1_CGC34_0_Prop8_0, in4526, M5_UM5_1_CC_1_CGC34_0_CGC23_line3);
or5 M5_UM5_1_CC_1_CGC34_0_CGC23_Ao5a_4(M5_UM5_1_CC_1_CGC34_0_LocalCarry33_27, M5_UM5_1_CC_1_CGC34_0_CGC23_line0, M5_UM5_1_CC_1_CGC34_0_CGC23_line1, M5_UM5_1_CC_1_CGC34_0_CGC23_line2, M5_UM5_1_CC_1_CGC34_0_CGC23_line3, CarryXbus_33);
and2 M5_UM5_1_CC_1_CGC34_1_CB5_0_Ao2_0(PropXbus_0, in4526, M5_UM5_1_CC_1_CGC34_1_CB5_0_line0);
or2 M5_UM5_1_CC_1_CGC34_1_CB5_0_Ao2_1(M5_GenXbus_0, M5_UM5_1_CC_1_CGC34_1_CB5_0_line0, CarryXbus_0);
and2 M5_UM5_1_CC_1_CGC34_1_CB5_1_Ao3a_0(PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_1_CGC34_1_CB5_1_line0);
and3 M5_UM5_1_CC_1_CGC34_1_CB5_1_Ao3a_1(PropXbus_1, PropXbus_0, in4526, M5_UM5_1_CC_1_CGC34_1_CB5_1_line1);
or3 M5_UM5_1_CC_1_CGC34_1_CB5_1_Ao3a_2(M5_GenXbus_1, M5_UM5_1_CC_1_CGC34_1_CB5_1_line0, M5_UM5_1_CC_1_CGC34_1_CB5_1_line1, CarryXbus_1);
and2 M5_UM5_1_CC_1_CGC34_1_CB5_2_Ao4a_0(PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_1_CGC34_1_CB5_2_line0);
and3 M5_UM5_1_CC_1_CGC34_1_CB5_2_Ao4a_1(PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_1_CGC34_1_CB5_2_line1);
and4 M5_UM5_1_CC_1_CGC34_1_CB5_2_Ao4a_2(PropXbus_2, PropXbus_1, PropXbus_0, in4526, M5_UM5_1_CC_1_CGC34_1_CB5_2_line2);
or4 M5_UM5_1_CC_1_CGC34_1_CB5_2_Ao4a_3(M5_GenXbus_2, M5_UM5_1_CC_1_CGC34_1_CB5_2_line0, M5_UM5_1_CC_1_CGC34_1_CB5_2_line1, M5_UM5_1_CC_1_CGC34_1_CB5_2_line2, CarryXbus_2);
and2 M5_UM5_1_CC_1_CGC34_1_CB5_3_Ao5a_0(PropXbus_3, M5_GenXbus_2, M5_UM5_1_CC_1_CGC34_1_CB5_3_line0);
and3 M5_UM5_1_CC_1_CGC34_1_CB5_3_Ao5a_1(PropXbus_3, PropXbus_2, M5_GenXbus_1, M5_UM5_1_CC_1_CGC34_1_CB5_3_line1);
and4 M5_UM5_1_CC_1_CGC34_1_CB5_3_Ao5a_2(PropXbus_3, PropXbus_2, PropXbus_1, M5_GenXbus_0, M5_UM5_1_CC_1_CGC34_1_CB5_3_line2);
and5 M5_UM5_1_CC_1_CGC34_1_CB5_3_Ao5a_3(PropXbus_3, PropXbus_2, PropXbus_1, PropXbus_0, in4526, M5_UM5_1_CC_1_CGC34_1_CB5_3_line3);
or5 M5_UM5_1_CC_1_CGC34_1_CB5_3_Ao5a_4(M5_GenXbus_3, M5_UM5_1_CC_1_CGC34_1_CB5_3_line0, M5_UM5_1_CC_1_CGC34_1_CB5_3_line1, M5_UM5_1_CC_1_CGC34_1_CB5_3_line2, M5_UM5_1_CC_1_CGC34_1_CB5_3_line3, CarryXbus_3);
and2 M5_UM5_1_CC_1_CGC34_2_CB5_0_Ao2_0(PropXbus_9, CarryXbus_8, M5_UM5_1_CC_1_CGC34_2_CB5_0_line0);
or2 M5_UM5_1_CC_1_CGC34_2_CB5_0_Ao2_1(M5_GenXbus_9, M5_UM5_1_CC_1_CGC34_2_CB5_0_line0, CarryXbus_9);
and2 M5_UM5_1_CC_1_CGC34_2_CB5_1_Ao3a_0(PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_1_CGC34_2_CB5_1_line0);
and3 M5_UM5_1_CC_1_CGC34_2_CB5_1_Ao3a_1(PropXbus_10, PropXbus_9, CarryXbus_8, M5_UM5_1_CC_1_CGC34_2_CB5_1_line1);
or3 M5_UM5_1_CC_1_CGC34_2_CB5_1_Ao3a_2(M5_GenXbus_10, M5_UM5_1_CC_1_CGC34_2_CB5_1_line0, M5_UM5_1_CC_1_CGC34_2_CB5_1_line1, CarryXbus_10);
and2 M5_UM5_1_CC_1_CGC34_2_CB5_2_Ao4a_0(PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_1_CGC34_2_CB5_2_line0);
and3 M5_UM5_1_CC_1_CGC34_2_CB5_2_Ao4a_1(PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_1_CGC34_2_CB5_2_line1);
and4 M5_UM5_1_CC_1_CGC34_2_CB5_2_Ao4a_2(PropXbus_11, PropXbus_10, PropXbus_9, CarryXbus_8, M5_UM5_1_CC_1_CGC34_2_CB5_2_line2);
or4 M5_UM5_1_CC_1_CGC34_2_CB5_2_Ao4a_3(M5_GenXbus_11, M5_UM5_1_CC_1_CGC34_2_CB5_2_line0, M5_UM5_1_CC_1_CGC34_2_CB5_2_line1, M5_UM5_1_CC_1_CGC34_2_CB5_2_line2, CarryXbus_11);
and2 M5_UM5_1_CC_1_CGC34_2_CB5_3_Ao5a_0(PropXbus_12, M5_GenXbus_11, M5_UM5_1_CC_1_CGC34_2_CB5_3_line0);
and3 M5_UM5_1_CC_1_CGC34_2_CB5_3_Ao5a_1(PropXbus_12, PropXbus_11, M5_GenXbus_10, M5_UM5_1_CC_1_CGC34_2_CB5_3_line1);
and4 M5_UM5_1_CC_1_CGC34_2_CB5_3_Ao5a_2(PropXbus_12, PropXbus_11, PropXbus_10, M5_GenXbus_9, M5_UM5_1_CC_1_CGC34_2_CB5_3_line2);
and5 M5_UM5_1_CC_1_CGC34_2_CB5_3_Ao5a_3(PropXbus_12, PropXbus_11, PropXbus_10, PropXbus_9, CarryXbus_8, M5_UM5_1_CC_1_CGC34_2_CB5_3_line3);
or5 M5_UM5_1_CC_1_CGC34_2_CB5_3_Ao5a_4(M5_GenXbus_12, M5_UM5_1_CC_1_CGC34_2_CB5_3_line0, M5_UM5_1_CC_1_CGC34_2_CB5_3_line1, M5_UM5_1_CC_1_CGC34_2_CB5_3_line2, M5_UM5_1_CC_1_CGC34_2_CB5_3_line3, CarryXbus_12);
and2 M5_UM5_1_CC_1_CGC34_3_CB5_0_Ao2_0(PropXbus_18, CarryXbus_17, M5_UM5_1_CC_1_CGC34_3_CB5_0_line0);
or2 M5_UM5_1_CC_1_CGC34_3_CB5_0_Ao2_1(M5_GenXbus_18, M5_UM5_1_CC_1_CGC34_3_CB5_0_line0, CarryXbus_18);
and2 M5_UM5_1_CC_1_CGC34_3_CB5_1_Ao3a_0(PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_1_CGC34_3_CB5_1_line0);
and3 M5_UM5_1_CC_1_CGC34_3_CB5_1_Ao3a_1(PropXbus_19, PropXbus_18, CarryXbus_17, M5_UM5_1_CC_1_CGC34_3_CB5_1_line1);
or3 M5_UM5_1_CC_1_CGC34_3_CB5_1_Ao3a_2(M5_GenXbus_19, M5_UM5_1_CC_1_CGC34_3_CB5_1_line0, M5_UM5_1_CC_1_CGC34_3_CB5_1_line1, CarryXbus_19);
and2 M5_UM5_1_CC_1_CGC34_3_CB5_2_Ao4a_0(PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_1_CGC34_3_CB5_2_line0);
and3 M5_UM5_1_CC_1_CGC34_3_CB5_2_Ao4a_1(PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_1_CGC34_3_CB5_2_line1);
and4 M5_UM5_1_CC_1_CGC34_3_CB5_2_Ao4a_2(PropXbus_20, PropXbus_19, PropXbus_18, CarryXbus_17, M5_UM5_1_CC_1_CGC34_3_CB5_2_line2);
or4 M5_UM5_1_CC_1_CGC34_3_CB5_2_Ao4a_3(M5_GenXbus_20, M5_UM5_1_CC_1_CGC34_3_CB5_2_line0, M5_UM5_1_CC_1_CGC34_3_CB5_2_line1, M5_UM5_1_CC_1_CGC34_3_CB5_2_line2, CarryXbus_20);
and2 M5_UM5_1_CC_1_CGC34_3_CB5_3_Ao5a_0(PropXbus_21, M5_GenXbus_20, M5_UM5_1_CC_1_CGC34_3_CB5_3_line0);
and3 M5_UM5_1_CC_1_CGC34_3_CB5_3_Ao5a_1(PropXbus_21, PropXbus_20, M5_GenXbus_19, M5_UM5_1_CC_1_CGC34_3_CB5_3_line1);
and4 M5_UM5_1_CC_1_CGC34_3_CB5_3_Ao5a_2(PropXbus_21, PropXbus_20, PropXbus_19, M5_GenXbus_18, M5_UM5_1_CC_1_CGC34_3_CB5_3_line2);
and5 M5_UM5_1_CC_1_CGC34_3_CB5_3_Ao5a_3(PropXbus_21, PropXbus_20, PropXbus_19, PropXbus_18, CarryXbus_17, M5_UM5_1_CC_1_CGC34_3_CB5_3_line3);
or5 M5_UM5_1_CC_1_CGC34_3_CB5_3_Ao5a_4(M5_GenXbus_21, M5_UM5_1_CC_1_CGC34_3_CB5_3_line0, M5_UM5_1_CC_1_CGC34_3_CB5_3_line1, M5_UM5_1_CC_1_CGC34_3_CB5_3_line2, M5_UM5_1_CC_1_CGC34_3_CB5_3_line3, CarryXbus_21);
and2 M5_UM5_1_CC_1_CGC34_4_CB5_0_Ao2_0(PropXbus_27, CarryXbus_26, M5_UM5_1_CC_1_CGC34_4_CB5_0_line0);
or2 M5_UM5_1_CC_1_CGC34_4_CB5_0_Ao2_1(M5_GenXbus_27, M5_UM5_1_CC_1_CGC34_4_CB5_0_line0, CarryXbus_27);
and2 M5_UM5_1_CC_1_CGC34_4_CB5_1_Ao3a_0(PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_1_CGC34_4_CB5_1_line0);
and3 M5_UM5_1_CC_1_CGC34_4_CB5_1_Ao3a_1(PropXbus_28, PropXbus_27, CarryXbus_26, M5_UM5_1_CC_1_CGC34_4_CB5_1_line1);
or3 M5_UM5_1_CC_1_CGC34_4_CB5_1_Ao3a_2(M5_GenXbus_28, M5_UM5_1_CC_1_CGC34_4_CB5_1_line0, M5_UM5_1_CC_1_CGC34_4_CB5_1_line1, CarryXbus_28);
and2 M5_UM5_1_CC_1_CGC34_4_CB5_2_Ao4a_0(PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_1_CGC34_4_CB5_2_line0);
and3 M5_UM5_1_CC_1_CGC34_4_CB5_2_Ao4a_1(PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_1_CGC34_4_CB5_2_line1);
and4 M5_UM5_1_CC_1_CGC34_4_CB5_2_Ao4a_2(PropXbus_29, PropXbus_28, PropXbus_27, CarryXbus_26, M5_UM5_1_CC_1_CGC34_4_CB5_2_line2);
or4 M5_UM5_1_CC_1_CGC34_4_CB5_2_Ao4a_3(M5_GenXbus_29, M5_UM5_1_CC_1_CGC34_4_CB5_2_line0, M5_UM5_1_CC_1_CGC34_4_CB5_2_line1, M5_UM5_1_CC_1_CGC34_4_CB5_2_line2, CarryXbus_29);
and2 M5_UM5_1_CC_1_CGC34_4_CB5_3_Ao5a_0(PropXbus_30, M5_GenXbus_29, M5_UM5_1_CC_1_CGC34_4_CB5_3_line0);
and3 M5_UM5_1_CC_1_CGC34_4_CB5_3_Ao5a_1(PropXbus_30, PropXbus_29, M5_GenXbus_28, M5_UM5_1_CC_1_CGC34_4_CB5_3_line1);
and4 M5_UM5_1_CC_1_CGC34_4_CB5_3_Ao5a_2(PropXbus_30, PropXbus_29, PropXbus_28, M5_GenXbus_27, M5_UM5_1_CC_1_CGC34_4_CB5_3_line2);
and5 M5_UM5_1_CC_1_CGC34_4_CB5_3_Ao5a_3(PropXbus_30, PropXbus_29, PropXbus_28, PropXbus_27, CarryXbus_26, M5_UM5_1_CC_1_CGC34_4_CB5_3_line3);
or5 M5_UM5_1_CC_1_CGC34_4_CB5_3_Ao5a_4(M5_GenXbus_30, M5_UM5_1_CC_1_CGC34_4_CB5_3_line0, M5_UM5_1_CC_1_CGC34_4_CB5_3_line1, M5_UM5_1_CC_1_CGC34_4_CB5_3_line2, M5_UM5_1_CC_1_CGC34_4_CB5_3_line3, CarryXbus_30);
inv M5_UM5_1_CC_2_Mux0(CarryXbus_31, M5_UM5_1_CC_2_Not_ContIn);
and2 M5_UM5_1_CC_2_Mux1(LocalCarryXCin0_33, M5_UM5_1_CC_2_Not_ContIn, M5_UM5_1_CC_2_line1);
and2 M5_UM5_1_CC_2_Mux2(LocalCarryXCin1_33, CarryXbus_31, M5_UM5_1_CC_2_line2);
or2 M5_UM5_1_CC_2_Mux3(M5_UM5_1_CC_2_line1, M5_UM5_1_CC_2_line2, out273);
inv M6_UM6_0_CSX6_0_Xo0(PropXbus_0, M6_UM6_0_CSX6_0_NotA);
inv M6_UM6_0_CSX6_0_Xo1(in4526, M6_UM6_0_CSX6_0_NotB);
nand2 M6_UM6_0_CSX6_0_Xo2(M6_UM6_0_CSX6_0_NotA, in4526, M6_UM6_0_CSX6_0_line2);
nand2 M6_UM6_0_CSX6_0_Xo3(M6_UM6_0_CSX6_0_NotB, PropXbus_0, M6_UM6_0_CSX6_0_line3);
nand2 M6_UM6_0_CSX6_0_Xo4(M6_UM6_0_CSX6_0_line2, M6_UM6_0_CSX6_0_line3, out373);
inv M6_UM6_0_CSX6_1_Xo0(PropXbus_1, M6_UM6_0_CSX6_1_NotA);
inv M6_UM6_0_CSX6_1_Xo1(CarryXbus_0, M6_UM6_0_CSX6_1_NotB);
nand2 M6_UM6_0_CSX6_1_Xo2(M6_UM6_0_CSX6_1_NotA, CarryXbus_0, M6_UM6_0_CSX6_1_line2);
nand2 M6_UM6_0_CSX6_1_Xo3(M6_UM6_0_CSX6_1_NotB, PropXbus_1, M6_UM6_0_CSX6_1_line3);
nand2 M6_UM6_0_CSX6_1_Xo4(M6_UM6_0_CSX6_1_line2, M6_UM6_0_CSX6_1_line3, out397);
inv M6_UM6_0_CSX6_2_Xo0(PropXbus_2, M6_UM6_0_CSX6_2_NotA);
inv M6_UM6_0_CSX6_2_Xo1(CarryXbus_1, M6_UM6_0_CSX6_2_NotB);
nand2 M6_UM6_0_CSX6_2_Xo2(M6_UM6_0_CSX6_2_NotA, CarryXbus_1, M6_UM6_0_CSX6_2_line2);
nand2 M6_UM6_0_CSX6_2_Xo3(M6_UM6_0_CSX6_2_NotB, PropXbus_2, M6_UM6_0_CSX6_2_line3);
nand2 M6_UM6_0_CSX6_2_Xo4(M6_UM6_0_CSX6_2_line2, M6_UM6_0_CSX6_2_line3, out394);
inv M6_UM6_0_CSX6_3_Xo0(PropXbus_3, M6_UM6_0_CSX6_3_NotA);
inv M6_UM6_0_CSX6_3_Xo1(CarryXbus_2, M6_UM6_0_CSX6_3_NotB);
nand2 M6_UM6_0_CSX6_3_Xo2(M6_UM6_0_CSX6_3_NotA, CarryXbus_2, M6_UM6_0_CSX6_3_line2);
nand2 M6_UM6_0_CSX6_3_Xo3(M6_UM6_0_CSX6_3_NotB, PropXbus_3, M6_UM6_0_CSX6_3_line3);
nand2 M6_UM6_0_CSX6_3_Xo4(M6_UM6_0_CSX6_3_line2, M6_UM6_0_CSX6_3_line3, out391);
inv M6_UM6_0_CSX6_4_Xo0(PropXbus_4, M6_UM6_0_CSX6_4_NotA);
inv M6_UM6_0_CSX6_4_Xo1(CarryXbus_3, M6_UM6_0_CSX6_4_NotB);
nand2 M6_UM6_0_CSX6_4_Xo2(M6_UM6_0_CSX6_4_NotA, CarryXbus_3, M6_UM6_0_CSX6_4_line2);
nand2 M6_UM6_0_CSX6_4_Xo3(M6_UM6_0_CSX6_4_NotB, PropXbus_4, M6_UM6_0_CSX6_4_line3);
nand2 M6_UM6_0_CSX6_4_Xo4(M6_UM6_0_CSX6_4_line2, M6_UM6_0_CSX6_4_line3, out388);
inv M6_UM6_0_CSX6_5_Xo0(PropXbus_5, M6_UM6_0_CSX6_5_NotA);
inv M6_UM6_0_CSX6_5_Xo1(CarryXbus_4, M6_UM6_0_CSX6_5_NotB);
nand2 M6_UM6_0_CSX6_5_Xo2(M6_UM6_0_CSX6_5_NotA, CarryXbus_4, M6_UM6_0_CSX6_5_line2);
nand2 M6_UM6_0_CSX6_5_Xo3(M6_UM6_0_CSX6_5_NotB, PropXbus_5, M6_UM6_0_CSX6_5_line3);
nand2 M6_UM6_0_CSX6_5_Xo4(M6_UM6_0_CSX6_5_line2, M6_UM6_0_CSX6_5_line3, out385);
inv M6_UM6_1_CSM4_0_Xo0(PropXbus_6, M6_UM6_1_CSM4_0_NotA);
inv M6_UM6_1_CSM4_0_Xo1(M5_GenXbus_5, M6_UM6_1_CSM4_0_NotB);
nand2 M6_UM6_1_CSM4_0_Xo2(M6_UM6_1_CSM4_0_NotA, M5_GenXbus_5, M6_UM6_1_CSM4_0_line2);
nand2 M6_UM6_1_CSM4_0_Xo3(M6_UM6_1_CSM4_0_NotB, PropXbus_6, M6_UM6_1_CSM4_0_line3);
nand2 M6_UM6_1_CSM4_0_Xo4(M6_UM6_1_CSM4_0_line2, M6_UM6_1_CSM4_0_line3, M6_UM6_1_Sum0_0);
inv M6_UM6_1_CSM4_1_Xo0(PropXbus_7, M6_UM6_1_CSM4_1_NotA);
inv M6_UM6_1_CSM4_1_Xo1(LocalCarryXCin0_6, M6_UM6_1_CSM4_1_NotB);
nand2 M6_UM6_1_CSM4_1_Xo2(M6_UM6_1_CSM4_1_NotA, LocalCarryXCin0_6, M6_UM6_1_CSM4_1_line2);
nand2 M6_UM6_1_CSM4_1_Xo3(M6_UM6_1_CSM4_1_NotB, PropXbus_7, M6_UM6_1_CSM4_1_line3);
nand2 M6_UM6_1_CSM4_1_Xo4(M6_UM6_1_CSM4_1_line2, M6_UM6_1_CSM4_1_line3, M6_UM6_1_Sum0_1);
inv M6_UM6_1_CSM4_2_Xo0(PropXbus_8, M6_UM6_1_CSM4_2_NotA);
inv M6_UM6_1_CSM4_2_Xo1(LocalCarryXCin0_7, M6_UM6_1_CSM4_2_NotB);
nand2 M6_UM6_1_CSM4_2_Xo2(M6_UM6_1_CSM4_2_NotA, LocalCarryXCin0_7, M6_UM6_1_CSM4_2_line2);
nand2 M6_UM6_1_CSM4_2_Xo3(M6_UM6_1_CSM4_2_NotB, PropXbus_8, M6_UM6_1_CSM4_2_line3);
nand2 M6_UM6_1_CSM4_2_Xo4(M6_UM6_1_CSM4_2_line2, M6_UM6_1_CSM4_2_line3, M6_UM6_1_Sum0_2);
inv M6_UM6_1_CSM4_3_Xo0(PropXbus_6, M6_UM6_1_CSM4_3_NotA);
inv M6_UM6_1_CSM4_3_Xo1(LocalCarryXCin1_5, M6_UM6_1_CSM4_3_NotB);
nand2 M6_UM6_1_CSM4_3_Xo2(M6_UM6_1_CSM4_3_NotA, LocalCarryXCin1_5, M6_UM6_1_CSM4_3_line2);
nand2 M6_UM6_1_CSM4_3_Xo3(M6_UM6_1_CSM4_3_NotB, PropXbus_6, M6_UM6_1_CSM4_3_line3);
nand2 M6_UM6_1_CSM4_3_Xo4(M6_UM6_1_CSM4_3_line2, M6_UM6_1_CSM4_3_line3, M6_UM6_1_Sum1_0);
inv M6_UM6_1_CSM4_4_Xo0(PropXbus_7, M6_UM6_1_CSM4_4_NotA);
inv M6_UM6_1_CSM4_4_Xo1(LocalCarryXCin1_6, M6_UM6_1_CSM4_4_NotB);
nand2 M6_UM6_1_CSM4_4_Xo2(M6_UM6_1_CSM4_4_NotA, LocalCarryXCin1_6, M6_UM6_1_CSM4_4_line2);
nand2 M6_UM6_1_CSM4_4_Xo3(M6_UM6_1_CSM4_4_NotB, PropXbus_7, M6_UM6_1_CSM4_4_line3);
nand2 M6_UM6_1_CSM4_4_Xo4(M6_UM6_1_CSM4_4_line2, M6_UM6_1_CSM4_4_line3, M6_UM6_1_Sum1_1);
inv M6_UM6_1_CSM4_5_Xo0(PropXbus_8, M6_UM6_1_CSM4_5_NotA);
inv M6_UM6_1_CSM4_5_Xo1(LocalCarryXCin1_7, M6_UM6_1_CSM4_5_NotB);
nand2 M6_UM6_1_CSM4_5_Xo2(M6_UM6_1_CSM4_5_NotA, LocalCarryXCin1_7, M6_UM6_1_CSM4_5_line2);
nand2 M6_UM6_1_CSM4_5_Xo3(M6_UM6_1_CSM4_5_NotB, PropXbus_8, M6_UM6_1_CSM4_5_line3);
nand2 M6_UM6_1_CSM4_5_Xo4(M6_UM6_1_CSM4_5_line2, M6_UM6_1_CSM4_5_line3, M6_UM6_1_Sum1_2);
inv M6_UM6_1_CSM4_6_Mux0(CarryXbus_4, M6_UM6_1_CSM4_6_Not_ContIn);
and2 M6_UM6_1_CSM4_6_Mux1(M6_UM6_1_Sum0_0, M6_UM6_1_CSM4_6_Not_ContIn, M6_UM6_1_CSM4_6_line1);
and2 M6_UM6_1_CSM4_6_Mux2(M6_UM6_1_Sum1_0, CarryXbus_4, M6_UM6_1_CSM4_6_line2);
or2 M6_UM6_1_CSM4_6_Mux3(M6_UM6_1_CSM4_6_line1, M6_UM6_1_CSM4_6_line2, out382);
inv M6_UM6_1_CSM4_7_Mux0(CarryXbus_4, M6_UM6_1_CSM4_7_Not_ContIn);
and2 M6_UM6_1_CSM4_7_Mux1(M6_UM6_1_Sum0_1, M6_UM6_1_CSM4_7_Not_ContIn, M6_UM6_1_CSM4_7_line1);
and2 M6_UM6_1_CSM4_7_Mux2(M6_UM6_1_Sum1_1, CarryXbus_4, M6_UM6_1_CSM4_7_line2);
or2 M6_UM6_1_CSM4_7_Mux3(M6_UM6_1_CSM4_7_line1, M6_UM6_1_CSM4_7_line2, out379);
inv M6_UM6_1_CSM4_8_Mux0(CarryXbus_4, M6_UM6_1_CSM4_8_Not_ContIn);
and2 M6_UM6_1_CSM4_8_Mux1(M6_UM6_1_Sum0_2, M6_UM6_1_CSM4_8_Not_ContIn, M6_UM6_1_CSM4_8_line1);
and2 M6_UM6_1_CSM4_8_Mux2(M6_UM6_1_Sum1_2, CarryXbus_4, M6_UM6_1_CSM4_8_line2);
or2 M6_UM6_1_CSM4_8_Mux3(M6_UM6_1_CSM4_8_line1, M6_UM6_1_CSM4_8_line2, out376);
inv M6_UM6_2_CSX6_0_Xo0(PropXbus_9, M6_UM6_2_CSX6_0_NotA);
inv M6_UM6_2_CSX6_0_Xo1(CarryXbus_8, M6_UM6_2_CSX6_0_NotB);
nand2 M6_UM6_2_CSX6_0_Xo2(M6_UM6_2_CSX6_0_NotA, CarryXbus_8, M6_UM6_2_CSX6_0_line2);
nand2 M6_UM6_2_CSX6_0_Xo3(M6_UM6_2_CSX6_0_NotB, PropXbus_9, M6_UM6_2_CSX6_0_line3);
nand2 M6_UM6_2_CSX6_0_Xo4(M6_UM6_2_CSX6_0_line2, M6_UM6_2_CSX6_0_line3, out344);
inv M6_UM6_2_CSX6_1_Xo0(PropXbus_10, M6_UM6_2_CSX6_1_NotA);
inv M6_UM6_2_CSX6_1_Xo1(CarryXbus_9, M6_UM6_2_CSX6_1_NotB);
nand2 M6_UM6_2_CSX6_1_Xo2(M6_UM6_2_CSX6_1_NotA, CarryXbus_9, M6_UM6_2_CSX6_1_line2);
nand2 M6_UM6_2_CSX6_1_Xo3(M6_UM6_2_CSX6_1_NotB, PropXbus_10, M6_UM6_2_CSX6_1_line3);
nand2 M6_UM6_2_CSX6_1_Xo4(M6_UM6_2_CSX6_1_line2, M6_UM6_2_CSX6_1_line3, out368);
inv M6_UM6_2_CSX6_2_Xo0(PropXbus_11, M6_UM6_2_CSX6_2_NotA);
inv M6_UM6_2_CSX6_2_Xo1(CarryXbus_10, M6_UM6_2_CSX6_2_NotB);
nand2 M6_UM6_2_CSX6_2_Xo2(M6_UM6_2_CSX6_2_NotA, CarryXbus_10, M6_UM6_2_CSX6_2_line2);
nand2 M6_UM6_2_CSX6_2_Xo3(M6_UM6_2_CSX6_2_NotB, PropXbus_11, M6_UM6_2_CSX6_2_line3);
nand2 M6_UM6_2_CSX6_2_Xo4(M6_UM6_2_CSX6_2_line2, M6_UM6_2_CSX6_2_line3, out365);
inv M6_UM6_2_CSX6_3_Xo0(PropXbus_12, M6_UM6_2_CSX6_3_NotA);
inv M6_UM6_2_CSX6_3_Xo1(CarryXbus_11, M6_UM6_2_CSX6_3_NotB);
nand2 M6_UM6_2_CSX6_3_Xo2(M6_UM6_2_CSX6_3_NotA, CarryXbus_11, M6_UM6_2_CSX6_3_line2);
nand2 M6_UM6_2_CSX6_3_Xo3(M6_UM6_2_CSX6_3_NotB, PropXbus_12, M6_UM6_2_CSX6_3_line3);
nand2 M6_UM6_2_CSX6_3_Xo4(M6_UM6_2_CSX6_3_line2, M6_UM6_2_CSX6_3_line3, out362);
inv M6_UM6_2_CSX6_4_Xo0(PropXbus_13, M6_UM6_2_CSX6_4_NotA);
inv M6_UM6_2_CSX6_4_Xo1(CarryXbus_12, M6_UM6_2_CSX6_4_NotB);
nand2 M6_UM6_2_CSX6_4_Xo2(M6_UM6_2_CSX6_4_NotA, CarryXbus_12, M6_UM6_2_CSX6_4_line2);
nand2 M6_UM6_2_CSX6_4_Xo3(M6_UM6_2_CSX6_4_NotB, PropXbus_13, M6_UM6_2_CSX6_4_line3);
nand2 M6_UM6_2_CSX6_4_Xo4(M6_UM6_2_CSX6_4_line2, M6_UM6_2_CSX6_4_line3, out359);
inv M6_UM6_2_CSX6_5_Xo0(PropXbus_14, M6_UM6_2_CSX6_5_NotA);
inv M6_UM6_2_CSX6_5_Xo1(CarryXbus_13, M6_UM6_2_CSX6_5_NotB);
nand2 M6_UM6_2_CSX6_5_Xo2(M6_UM6_2_CSX6_5_NotA, CarryXbus_13, M6_UM6_2_CSX6_5_line2);
nand2 M6_UM6_2_CSX6_5_Xo3(M6_UM6_2_CSX6_5_NotB, PropXbus_14, M6_UM6_2_CSX6_5_line3);
nand2 M6_UM6_2_CSX6_5_Xo4(M6_UM6_2_CSX6_5_line2, M6_UM6_2_CSX6_5_line3, out356);
inv M6_UM6_3_CSM4_0_Xo0(PropXbus_15, M6_UM6_3_CSM4_0_NotA);
inv M6_UM6_3_CSM4_0_Xo1(M5_GenXbus_14, M6_UM6_3_CSM4_0_NotB);
nand2 M6_UM6_3_CSM4_0_Xo2(M6_UM6_3_CSM4_0_NotA, M5_GenXbus_14, M6_UM6_3_CSM4_0_line2);
nand2 M6_UM6_3_CSM4_0_Xo3(M6_UM6_3_CSM4_0_NotB, PropXbus_15, M6_UM6_3_CSM4_0_line3);
nand2 M6_UM6_3_CSM4_0_Xo4(M6_UM6_3_CSM4_0_line2, M6_UM6_3_CSM4_0_line3, M6_UM6_3_Sum0_0);
inv M6_UM6_3_CSM4_1_Xo0(PropXbus_16, M6_UM6_3_CSM4_1_NotA);
inv M6_UM6_3_CSM4_1_Xo1(LocalCarryXCin0_15, M6_UM6_3_CSM4_1_NotB);
nand2 M6_UM6_3_CSM4_1_Xo2(M6_UM6_3_CSM4_1_NotA, LocalCarryXCin0_15, M6_UM6_3_CSM4_1_line2);
nand2 M6_UM6_3_CSM4_1_Xo3(M6_UM6_3_CSM4_1_NotB, PropXbus_16, M6_UM6_3_CSM4_1_line3);
nand2 M6_UM6_3_CSM4_1_Xo4(M6_UM6_3_CSM4_1_line2, M6_UM6_3_CSM4_1_line3, M6_UM6_3_Sum0_1);
inv M6_UM6_3_CSM4_2_Xo0(PropXbus_17, M6_UM6_3_CSM4_2_NotA);
inv M6_UM6_3_CSM4_2_Xo1(LocalCarryXCin0_16, M6_UM6_3_CSM4_2_NotB);
nand2 M6_UM6_3_CSM4_2_Xo2(M6_UM6_3_CSM4_2_NotA, LocalCarryXCin0_16, M6_UM6_3_CSM4_2_line2);
nand2 M6_UM6_3_CSM4_2_Xo3(M6_UM6_3_CSM4_2_NotB, PropXbus_17, M6_UM6_3_CSM4_2_line3);
nand2 M6_UM6_3_CSM4_2_Xo4(M6_UM6_3_CSM4_2_line2, M6_UM6_3_CSM4_2_line3, M6_UM6_3_Sum0_2);
inv M6_UM6_3_CSM4_3_Xo0(PropXbus_15, M6_UM6_3_CSM4_3_NotA);
inv M6_UM6_3_CSM4_3_Xo1(LocalCarryXCin1_14, M6_UM6_3_CSM4_3_NotB);
nand2 M6_UM6_3_CSM4_3_Xo2(M6_UM6_3_CSM4_3_NotA, LocalCarryXCin1_14, M6_UM6_3_CSM4_3_line2);
nand2 M6_UM6_3_CSM4_3_Xo3(M6_UM6_3_CSM4_3_NotB, PropXbus_15, M6_UM6_3_CSM4_3_line3);
nand2 M6_UM6_3_CSM4_3_Xo4(M6_UM6_3_CSM4_3_line2, M6_UM6_3_CSM4_3_line3, M6_UM6_3_Sum1_0);
inv M6_UM6_3_CSM4_4_Xo0(PropXbus_16, M6_UM6_3_CSM4_4_NotA);
inv M6_UM6_3_CSM4_4_Xo1(LocalCarryXCin1_15, M6_UM6_3_CSM4_4_NotB);
nand2 M6_UM6_3_CSM4_4_Xo2(M6_UM6_3_CSM4_4_NotA, LocalCarryXCin1_15, M6_UM6_3_CSM4_4_line2);
nand2 M6_UM6_3_CSM4_4_Xo3(M6_UM6_3_CSM4_4_NotB, PropXbus_16, M6_UM6_3_CSM4_4_line3);
nand2 M6_UM6_3_CSM4_4_Xo4(M6_UM6_3_CSM4_4_line2, M6_UM6_3_CSM4_4_line3, M6_UM6_3_Sum1_1);
inv M6_UM6_3_CSM4_5_Xo0(PropXbus_17, M6_UM6_3_CSM4_5_NotA);
inv M6_UM6_3_CSM4_5_Xo1(LocalCarryXCin1_16, M6_UM6_3_CSM4_5_NotB);
nand2 M6_UM6_3_CSM4_5_Xo2(M6_UM6_3_CSM4_5_NotA, LocalCarryXCin1_16, M6_UM6_3_CSM4_5_line2);
nand2 M6_UM6_3_CSM4_5_Xo3(M6_UM6_3_CSM4_5_NotB, PropXbus_17, M6_UM6_3_CSM4_5_line3);
nand2 M6_UM6_3_CSM4_5_Xo4(M6_UM6_3_CSM4_5_line2, M6_UM6_3_CSM4_5_line3, M6_UM6_3_Sum1_2);
inv M6_UM6_3_CSM4_6_Mux0(CarryXbus_13, M6_UM6_3_CSM4_6_Not_ContIn);
and2 M6_UM6_3_CSM4_6_Mux1(M6_UM6_3_Sum0_0, M6_UM6_3_CSM4_6_Not_ContIn, M6_UM6_3_CSM4_6_line1);
and2 M6_UM6_3_CSM4_6_Mux2(M6_UM6_3_Sum1_0, CarryXbus_13, M6_UM6_3_CSM4_6_line2);
or2 M6_UM6_3_CSM4_6_Mux3(M6_UM6_3_CSM4_6_line1, M6_UM6_3_CSM4_6_line2, out353);
inv M6_UM6_3_CSM4_7_Mux0(CarryXbus_13, M6_UM6_3_CSM4_7_Not_ContIn);
and2 M6_UM6_3_CSM4_7_Mux1(M6_UM6_3_Sum0_1, M6_UM6_3_CSM4_7_Not_ContIn, M6_UM6_3_CSM4_7_line1);
and2 M6_UM6_3_CSM4_7_Mux2(M6_UM6_3_Sum1_1, CarryXbus_13, M6_UM6_3_CSM4_7_line2);
or2 M6_UM6_3_CSM4_7_Mux3(M6_UM6_3_CSM4_7_line1, M6_UM6_3_CSM4_7_line2, out350);
inv M6_UM6_3_CSM4_8_Mux0(CarryXbus_13, M6_UM6_3_CSM4_8_Not_ContIn);
and2 M6_UM6_3_CSM4_8_Mux1(M6_UM6_3_Sum0_2, M6_UM6_3_CSM4_8_Not_ContIn, M6_UM6_3_CSM4_8_line1);
and2 M6_UM6_3_CSM4_8_Mux2(M6_UM6_3_Sum1_2, CarryXbus_13, M6_UM6_3_CSM4_8_line2);
or2 M6_UM6_3_CSM4_8_Mux3(M6_UM6_3_CSM4_8_line1, M6_UM6_3_CSM4_8_line2, out347);
inv M6_UM6_4_CSX6_0_Xo0(PropXbus_18, M6_UM6_4_CSX6_0_NotA);
inv M6_UM6_4_CSX6_0_Xo1(CarryXbus_17, M6_UM6_4_CSX6_0_NotB);
nand2 M6_UM6_4_CSX6_0_Xo2(M6_UM6_4_CSX6_0_NotA, CarryXbus_17, M6_UM6_4_CSX6_0_line2);
nand2 M6_UM6_4_CSX6_0_Xo3(M6_UM6_4_CSX6_0_NotB, PropXbus_18, M6_UM6_4_CSX6_0_line3);
nand2 M6_UM6_4_CSX6_0_Xo4(M6_UM6_4_CSX6_0_line2, M6_UM6_4_CSX6_0_line3, out295);
inv M6_UM6_4_CSX6_1_Xo0(PropXbus_19, M6_UM6_4_CSX6_1_NotA);
inv M6_UM6_4_CSX6_1_Xo1(CarryXbus_18, M6_UM6_4_CSX6_1_NotB);
nand2 M6_UM6_4_CSX6_1_Xo2(M6_UM6_4_CSX6_1_NotA, CarryXbus_18, M6_UM6_4_CSX6_1_line2);
nand2 M6_UM6_4_CSX6_1_Xo3(M6_UM6_4_CSX6_1_NotB, PropXbus_19, M6_UM6_4_CSX6_1_line3);
nand2 M6_UM6_4_CSX6_1_Xo4(M6_UM6_4_CSX6_1_line2, M6_UM6_4_CSX6_1_line3, out319);
inv M6_UM6_4_CSX6_2_Xo0(PropXbus_20, M6_UM6_4_CSX6_2_NotA);
inv M6_UM6_4_CSX6_2_Xo1(CarryXbus_19, M6_UM6_4_CSX6_2_NotB);
nand2 M6_UM6_4_CSX6_2_Xo2(M6_UM6_4_CSX6_2_NotA, CarryXbus_19, M6_UM6_4_CSX6_2_line2);
nand2 M6_UM6_4_CSX6_2_Xo3(M6_UM6_4_CSX6_2_NotB, PropXbus_20, M6_UM6_4_CSX6_2_line3);
nand2 M6_UM6_4_CSX6_2_Xo4(M6_UM6_4_CSX6_2_line2, M6_UM6_4_CSX6_2_line3, out316);
inv M6_UM6_4_CSX6_3_Xo0(PropXbus_21, M6_UM6_4_CSX6_3_NotA);
inv M6_UM6_4_CSX6_3_Xo1(CarryXbus_20, M6_UM6_4_CSX6_3_NotB);
nand2 M6_UM6_4_CSX6_3_Xo2(M6_UM6_4_CSX6_3_NotA, CarryXbus_20, M6_UM6_4_CSX6_3_line2);
nand2 M6_UM6_4_CSX6_3_Xo3(M6_UM6_4_CSX6_3_NotB, PropXbus_21, M6_UM6_4_CSX6_3_line3);
nand2 M6_UM6_4_CSX6_3_Xo4(M6_UM6_4_CSX6_3_line2, M6_UM6_4_CSX6_3_line3, out313);
inv M6_UM6_4_CSX6_4_Xo0(PropXbus_22, M6_UM6_4_CSX6_4_NotA);
inv M6_UM6_4_CSX6_4_Xo1(CarryXbus_21, M6_UM6_4_CSX6_4_NotB);
nand2 M6_UM6_4_CSX6_4_Xo2(M6_UM6_4_CSX6_4_NotA, CarryXbus_21, M6_UM6_4_CSX6_4_line2);
nand2 M6_UM6_4_CSX6_4_Xo3(M6_UM6_4_CSX6_4_NotB, PropXbus_22, M6_UM6_4_CSX6_4_line3);
nand2 M6_UM6_4_CSX6_4_Xo4(M6_UM6_4_CSX6_4_line2, M6_UM6_4_CSX6_4_line3, out310);
inv M6_UM6_4_CSX6_5_Xo0(PropXbus_23, M6_UM6_4_CSX6_5_NotA);
inv M6_UM6_4_CSX6_5_Xo1(CarryXbus_22, M6_UM6_4_CSX6_5_NotB);
nand2 M6_UM6_4_CSX6_5_Xo2(M6_UM6_4_CSX6_5_NotA, CarryXbus_22, M6_UM6_4_CSX6_5_line2);
nand2 M6_UM6_4_CSX6_5_Xo3(M6_UM6_4_CSX6_5_NotB, PropXbus_23, M6_UM6_4_CSX6_5_line3);
nand2 M6_UM6_4_CSX6_5_Xo4(M6_UM6_4_CSX6_5_line2, M6_UM6_4_CSX6_5_line3, out307);
inv M6_UM6_5_CSM4_0_Xo0(PropXbus_24, M6_UM6_5_CSM4_0_NotA);
inv M6_UM6_5_CSM4_0_Xo1(M5_GenXbus_23, M6_UM6_5_CSM4_0_NotB);
nand2 M6_UM6_5_CSM4_0_Xo2(M6_UM6_5_CSM4_0_NotA, M5_GenXbus_23, M6_UM6_5_CSM4_0_line2);
nand2 M6_UM6_5_CSM4_0_Xo3(M6_UM6_5_CSM4_0_NotB, PropXbus_24, M6_UM6_5_CSM4_0_line3);
nand2 M6_UM6_5_CSM4_0_Xo4(M6_UM6_5_CSM4_0_line2, M6_UM6_5_CSM4_0_line3, M6_UM6_5_Sum0_0);
inv M6_UM6_5_CSM4_1_Xo0(PropXbus_25, M6_UM6_5_CSM4_1_NotA);
inv M6_UM6_5_CSM4_1_Xo1(LocalCarryXCin0_24, M6_UM6_5_CSM4_1_NotB);
nand2 M6_UM6_5_CSM4_1_Xo2(M6_UM6_5_CSM4_1_NotA, LocalCarryXCin0_24, M6_UM6_5_CSM4_1_line2);
nand2 M6_UM6_5_CSM4_1_Xo3(M6_UM6_5_CSM4_1_NotB, PropXbus_25, M6_UM6_5_CSM4_1_line3);
nand2 M6_UM6_5_CSM4_1_Xo4(M6_UM6_5_CSM4_1_line2, M6_UM6_5_CSM4_1_line3, M6_UM6_5_Sum0_1);
inv M6_UM6_5_CSM4_2_Xo0(PropXbus_26, M6_UM6_5_CSM4_2_NotA);
inv M6_UM6_5_CSM4_2_Xo1(LocalCarryXCin0_25, M6_UM6_5_CSM4_2_NotB);
nand2 M6_UM6_5_CSM4_2_Xo2(M6_UM6_5_CSM4_2_NotA, LocalCarryXCin0_25, M6_UM6_5_CSM4_2_line2);
nand2 M6_UM6_5_CSM4_2_Xo3(M6_UM6_5_CSM4_2_NotB, PropXbus_26, M6_UM6_5_CSM4_2_line3);
nand2 M6_UM6_5_CSM4_2_Xo4(M6_UM6_5_CSM4_2_line2, M6_UM6_5_CSM4_2_line3, M6_UM6_5_Sum0_2);
inv M6_UM6_5_CSM4_3_Xo0(PropXbus_24, M6_UM6_5_CSM4_3_NotA);
inv M6_UM6_5_CSM4_3_Xo1(LocalCarryXCin1_23, M6_UM6_5_CSM4_3_NotB);
nand2 M6_UM6_5_CSM4_3_Xo2(M6_UM6_5_CSM4_3_NotA, LocalCarryXCin1_23, M6_UM6_5_CSM4_3_line2);
nand2 M6_UM6_5_CSM4_3_Xo3(M6_UM6_5_CSM4_3_NotB, PropXbus_24, M6_UM6_5_CSM4_3_line3);
nand2 M6_UM6_5_CSM4_3_Xo4(M6_UM6_5_CSM4_3_line2, M6_UM6_5_CSM4_3_line3, M6_UM6_5_Sum1_0);
inv M6_UM6_5_CSM4_4_Xo0(PropXbus_25, M6_UM6_5_CSM4_4_NotA);
inv M6_UM6_5_CSM4_4_Xo1(LocalCarryXCin1_24, M6_UM6_5_CSM4_4_NotB);
nand2 M6_UM6_5_CSM4_4_Xo2(M6_UM6_5_CSM4_4_NotA, LocalCarryXCin1_24, M6_UM6_5_CSM4_4_line2);
nand2 M6_UM6_5_CSM4_4_Xo3(M6_UM6_5_CSM4_4_NotB, PropXbus_25, M6_UM6_5_CSM4_4_line3);
nand2 M6_UM6_5_CSM4_4_Xo4(M6_UM6_5_CSM4_4_line2, M6_UM6_5_CSM4_4_line3, M6_UM6_5_Sum1_1);
inv M6_UM6_5_CSM4_5_Xo0(PropXbus_26, M6_UM6_5_CSM4_5_NotA);
inv M6_UM6_5_CSM4_5_Xo1(LocalCarryXCin1_25, M6_UM6_5_CSM4_5_NotB);
nand2 M6_UM6_5_CSM4_5_Xo2(M6_UM6_5_CSM4_5_NotA, LocalCarryXCin1_25, M6_UM6_5_CSM4_5_line2);
nand2 M6_UM6_5_CSM4_5_Xo3(M6_UM6_5_CSM4_5_NotB, PropXbus_26, M6_UM6_5_CSM4_5_line3);
nand2 M6_UM6_5_CSM4_5_Xo4(M6_UM6_5_CSM4_5_line2, M6_UM6_5_CSM4_5_line3, M6_UM6_5_Sum1_2);
inv M6_UM6_5_CSM4_6_Mux0(CarryXbus_22, M6_UM6_5_CSM4_6_Not_ContIn);
and2 M6_UM6_5_CSM4_6_Mux1(M6_UM6_5_Sum0_0, M6_UM6_5_CSM4_6_Not_ContIn, M6_UM6_5_CSM4_6_line1);
and2 M6_UM6_5_CSM4_6_Mux2(M6_UM6_5_Sum1_0, CarryXbus_22, M6_UM6_5_CSM4_6_line2);
or2 M6_UM6_5_CSM4_6_Mux3(M6_UM6_5_CSM4_6_line1, M6_UM6_5_CSM4_6_line2, out304);
inv M6_UM6_5_CSM4_7_Mux0(CarryXbus_22, M6_UM6_5_CSM4_7_Not_ContIn);
and2 M6_UM6_5_CSM4_7_Mux1(M6_UM6_5_Sum0_1, M6_UM6_5_CSM4_7_Not_ContIn, M6_UM6_5_CSM4_7_line1);
and2 M6_UM6_5_CSM4_7_Mux2(M6_UM6_5_Sum1_1, CarryXbus_22, M6_UM6_5_CSM4_7_line2);
or2 M6_UM6_5_CSM4_7_Mux3(M6_UM6_5_CSM4_7_line1, M6_UM6_5_CSM4_7_line2, out301);
inv M6_UM6_5_CSM4_8_Mux0(CarryXbus_22, M6_UM6_5_CSM4_8_Not_ContIn);
and2 M6_UM6_5_CSM4_8_Mux1(M6_UM6_5_Sum0_2, M6_UM6_5_CSM4_8_Not_ContIn, M6_UM6_5_CSM4_8_line1);
and2 M6_UM6_5_CSM4_8_Mux2(M6_UM6_5_Sum1_2, CarryXbus_22, M6_UM6_5_CSM4_8_line2);
or2 M6_UM6_5_CSM4_8_Mux3(M6_UM6_5_CSM4_8_line1, M6_UM6_5_CSM4_8_line2, out298);
inv M6_UM6_6_CSX6_0_Xo0(PropXbus_27, M6_UM6_6_CSX6_0_NotA);
inv M6_UM6_6_CSX6_0_Xo1(CarryXbus_26, M6_UM6_6_CSX6_0_NotB);
nand2 M6_UM6_6_CSX6_0_Xo2(M6_UM6_6_CSX6_0_NotA, CarryXbus_26, M6_UM6_6_CSX6_0_line2);
nand2 M6_UM6_6_CSX6_0_Xo3(M6_UM6_6_CSX6_0_NotB, PropXbus_27, M6_UM6_6_CSX6_0_line3);
nand2 M6_UM6_6_CSX6_0_Xo4(M6_UM6_6_CSX6_0_line2, M6_UM6_6_CSX6_0_line3, out324);
inv M6_UM6_6_CSX6_1_Xo0(PropXbus_28, M6_UM6_6_CSX6_1_NotA);
inv M6_UM6_6_CSX6_1_Xo1(CarryXbus_27, M6_UM6_6_CSX6_1_NotB);
nand2 M6_UM6_6_CSX6_1_Xo2(M6_UM6_6_CSX6_1_NotA, CarryXbus_27, M6_UM6_6_CSX6_1_line2);
nand2 M6_UM6_6_CSX6_1_Xo3(M6_UM6_6_CSX6_1_NotB, PropXbus_28, M6_UM6_6_CSX6_1_line3);
nand2 M6_UM6_6_CSX6_1_Xo4(M6_UM6_6_CSX6_1_line2, M6_UM6_6_CSX6_1_line3, out336);
inv M6_UM6_6_CSX6_2_Xo0(PropXbus_29, M6_UM6_6_CSX6_2_NotA);
inv M6_UM6_6_CSX6_2_Xo1(CarryXbus_28, M6_UM6_6_CSX6_2_NotB);
nand2 M6_UM6_6_CSX6_2_Xo2(M6_UM6_6_CSX6_2_NotA, CarryXbus_28, M6_UM6_6_CSX6_2_line2);
nand2 M6_UM6_6_CSX6_2_Xo3(M6_UM6_6_CSX6_2_NotB, PropXbus_29, M6_UM6_6_CSX6_2_line3);
nand2 M6_UM6_6_CSX6_2_Xo4(M6_UM6_6_CSX6_2_line2, M6_UM6_6_CSX6_2_line3, out333);
inv M6_UM6_6_CSX6_3_Xo0(PropXbus_30, M6_UM6_6_CSX6_3_NotA);
inv M6_UM6_6_CSX6_3_Xo1(CarryXbus_29, M6_UM6_6_CSX6_3_NotB);
nand2 M6_UM6_6_CSX6_3_Xo2(M6_UM6_6_CSX6_3_NotA, CarryXbus_29, M6_UM6_6_CSX6_3_line2);
nand2 M6_UM6_6_CSX6_3_Xo3(M6_UM6_6_CSX6_3_NotB, PropXbus_30, M6_UM6_6_CSX6_3_line3);
nand2 M6_UM6_6_CSX6_3_Xo4(M6_UM6_6_CSX6_3_line2, M6_UM6_6_CSX6_3_line3, out330);
inv M6_UM6_6_CSX6_4_Xo0(PropXbus_31, M6_UM6_6_CSX6_4_NotA);
inv M6_UM6_6_CSX6_4_Xo1(CarryXbus_30, M6_UM6_6_CSX6_4_NotB);
nand2 M6_UM6_6_CSX6_4_Xo2(M6_UM6_6_CSX6_4_NotA, CarryXbus_30, M6_UM6_6_CSX6_4_line2);
nand2 M6_UM6_6_CSX6_4_Xo3(M6_UM6_6_CSX6_4_NotB, PropXbus_31, M6_UM6_6_CSX6_4_line3);
nand2 M6_UM6_6_CSX6_4_Xo4(M6_UM6_6_CSX6_4_line2, M6_UM6_6_CSX6_4_line3, out327);
inv M6_UM6_6_CSX6_5_Xo0(PropXbus_32, M6_UM6_6_CSX6_5_NotA);
inv M6_UM6_6_CSX6_5_Xo1(CarryXbus_31, M6_UM6_6_CSX6_5_NotB);
nand2 M6_UM6_6_CSX6_5_Xo2(M6_UM6_6_CSX6_5_NotA, CarryXbus_31, M6_UM6_6_CSX6_5_line2);
nand2 M6_UM6_6_CSX6_5_Xo3(M6_UM6_6_CSX6_5_NotB, PropXbus_32, M6_UM6_6_CSX6_5_line3);
nand2 M6_UM6_6_CSX6_5_Xo4(M6_UM6_6_CSX6_5_line2, M6_UM6_6_CSX6_5_line3, out471);
inv M6_UM6_7_Xo0(PropXbus_33, M6_UM6_7_NotA);
inv M6_UM6_7_Xo1(M5_GenXbus_32, M6_UM6_7_NotB);
nand2 M6_UM6_7_Xo2(M6_UM6_7_NotA, M5_GenXbus_32, M6_UM6_7_line2);
nand2 M6_UM6_7_Xo3(M6_UM6_7_NotB, PropXbus_33, M6_UM6_7_line3);
nand2 M6_UM6_7_Xo4(M6_UM6_7_line2, M6_UM6_7_line3, M6_Sum33_0);
inv M6_UM6_8_Xo0(PropXbus_33, M6_UM6_8_NotA);
inv M6_UM6_8_Xo1(LocalCarryXCin1_32, M6_UM6_8_NotB);
nand2 M6_UM6_8_Xo2(M6_UM6_8_NotA, LocalCarryXCin1_32, M6_UM6_8_line2);
nand2 M6_UM6_8_Xo3(M6_UM6_8_NotB, PropXbus_33, M6_UM6_8_line3);
nand2 M6_UM6_8_Xo4(M6_UM6_8_line2, M6_UM6_8_line3, M6_Sum33_1);
inv M6_UM6_9_Mux0(CarryXbus_31, M6_UM6_9_Not_ContIn);
and2 M6_UM6_9_Mux1(M6_Sum33_0, M6_UM6_9_Not_ContIn, M6_UM6_9_line1);
and2 M6_UM6_9_Mux2(M6_Sum33_1, CarryXbus_31, M6_UM6_9_line2);
or2 M6_UM6_9_Mux3(M6_UM6_9_line1, M6_UM6_9_line2, out469);
inv M7_GSP0_SP9nc0_SP7nc0_Xo0(M5_GenXbus_0, M7_GSP0_SP9nc0_SP7nc0_NotA);
inv M7_GSP0_SP9nc0_SP7nc0_Xo1(LocalCarryXCin0_1, M7_GSP0_SP9nc0_SP7nc0_NotB);
nand2 M7_GSP0_SP9nc0_SP7nc0_Xo2(M7_GSP0_SP9nc0_SP7nc0_NotA, LocalCarryXCin0_1, M7_GSP0_SP9nc0_SP7nc0_line2);
nand2 M7_GSP0_SP9nc0_SP7nc0_Xo3(M7_GSP0_SP9nc0_SP7nc0_NotB, M5_GenXbus_0, M7_GSP0_SP9nc0_SP7nc0_line3);
nand2 M7_GSP0_SP9nc0_SP7nc0_Xo4(M7_GSP0_SP9nc0_SP7nc0_line2, M7_GSP0_SP9nc0_SP7nc0_line3, M7_GSP0_SP9nc0_line0);
inv M7_GSP0_SP9nc0_SP7nc1_Xo0(LocalCarryXCin0_2, M7_GSP0_SP9nc0_SP7nc1_NotA);
inv M7_GSP0_SP9nc0_SP7nc1_Xo1(M7_GSP0_SP9nc0_line0, M7_GSP0_SP9nc0_SP7nc1_NotB);
nand2 M7_GSP0_SP9nc0_SP7nc1_Xo2(M7_GSP0_SP9nc0_SP7nc1_NotA, M7_GSP0_SP9nc0_line0, M7_GSP0_SP9nc0_SP7nc1_line2);
nand2 M7_GSP0_SP9nc0_SP7nc1_Xo3(M7_GSP0_SP9nc0_SP7nc1_NotB, LocalCarryXCin0_2, M7_GSP0_SP9nc0_SP7nc1_line3);
nand2 M7_GSP0_SP9nc0_SP7nc1_Xo4(M7_GSP0_SP9nc0_SP7nc1_line2, M7_GSP0_SP9nc0_SP7nc1_line3, M7_GSP0_SP9nc0_line1);
inv M7_GSP0_SP9nc0_SP7nc2_Xo0(LocalCarryXCin0_3, M7_GSP0_SP9nc0_SP7nc2_NotA);
inv M7_GSP0_SP9nc0_SP7nc2_Xo1(M7_GSP0_SP9nc0_line1, M7_GSP0_SP9nc0_SP7nc2_NotB);
nand2 M7_GSP0_SP9nc0_SP7nc2_Xo2(M7_GSP0_SP9nc0_SP7nc2_NotA, M7_GSP0_SP9nc0_line1, M7_GSP0_SP9nc0_SP7nc2_line2);
nand2 M7_GSP0_SP9nc0_SP7nc2_Xo3(M7_GSP0_SP9nc0_SP7nc2_NotB, LocalCarryXCin0_3, M7_GSP0_SP9nc0_SP7nc2_line3);
nand2 M7_GSP0_SP9nc0_SP7nc2_Xo4(M7_GSP0_SP9nc0_SP7nc2_line2, M7_GSP0_SP9nc0_SP7nc2_line3, M7_GSP0_SP9nc0_line2);
inv M7_GSP0_SP9nc0_SP7nc3_Xo0(PropXbus_0, M7_GSP0_SP9nc0_SP7nc3_NotA);
inv M7_GSP0_SP9nc0_SP7nc3_Xo1(M7_GSP0_SP9nc0_line2, M7_GSP0_SP9nc0_SP7nc3_NotB);
nand2 M7_GSP0_SP9nc0_SP7nc3_Xo2(M7_GSP0_SP9nc0_SP7nc3_NotA, M7_GSP0_SP9nc0_line2, M7_GSP0_SP9nc0_SP7nc3_line2);
nand2 M7_GSP0_SP9nc0_SP7nc3_Xo3(M7_GSP0_SP9nc0_SP7nc3_NotB, PropXbus_0, M7_GSP0_SP9nc0_SP7nc3_line3);
nand2 M7_GSP0_SP9nc0_SP7nc3_Xo4(M7_GSP0_SP9nc0_SP7nc3_line2, M7_GSP0_SP9nc0_SP7nc3_line3, M7_GSP0_SP9nc0_line3);
inv M7_GSP0_SP9nc0_SP7nc4_Xo0(PropXbus_1, M7_GSP0_SP9nc0_SP7nc4_NotA);
inv M7_GSP0_SP9nc0_SP7nc4_Xo1(M7_GSP0_SP9nc0_line3, M7_GSP0_SP9nc0_SP7nc4_NotB);
nand2 M7_GSP0_SP9nc0_SP7nc4_Xo2(M7_GSP0_SP9nc0_SP7nc4_NotA, M7_GSP0_SP9nc0_line3, M7_GSP0_SP9nc0_SP7nc4_line2);
nand2 M7_GSP0_SP9nc0_SP7nc4_Xo3(M7_GSP0_SP9nc0_SP7nc4_NotB, PropXbus_1, M7_GSP0_SP9nc0_SP7nc4_line3);
nand2 M7_GSP0_SP9nc0_SP7nc4_Xo4(M7_GSP0_SP9nc0_SP7nc4_line2, M7_GSP0_SP9nc0_SP7nc4_line3, M7_GSP0_SP9nc0_line4);
inv M7_GSP0_SP9nc0_SP7nc5_Xo0(PropXbus_2, M7_GSP0_SP9nc0_SP7nc5_NotA);
inv M7_GSP0_SP9nc0_SP7nc5_Xo1(M7_GSP0_SP9nc0_line4, M7_GSP0_SP9nc0_SP7nc5_NotB);
nand2 M7_GSP0_SP9nc0_SP7nc5_Xo2(M7_GSP0_SP9nc0_SP7nc5_NotA, M7_GSP0_SP9nc0_line4, M7_GSP0_SP9nc0_SP7nc5_line2);
nand2 M7_GSP0_SP9nc0_SP7nc5_Xo3(M7_GSP0_SP9nc0_SP7nc5_NotB, PropXbus_2, M7_GSP0_SP9nc0_SP7nc5_line3);
nand2 M7_GSP0_SP9nc0_SP7nc5_Xo4(M7_GSP0_SP9nc0_SP7nc5_line2, M7_GSP0_SP9nc0_SP7nc5_line3, M7_GSP0_line0);
inv M7_GSP0_SP9nc1_Xo0(PropXbus_3, M7_GSP0_SP9nc1_NotA);
inv M7_GSP0_SP9nc1_Xo1(M7_GSP0_line0, M7_GSP0_SP9nc1_NotB);
nand2 M7_GSP0_SP9nc1_Xo2(M7_GSP0_SP9nc1_NotA, M7_GSP0_line0, M7_GSP0_SP9nc1_line2);
nand2 M7_GSP0_SP9nc1_Xo3(M7_GSP0_SP9nc1_NotB, PropXbus_3, M7_GSP0_SP9nc1_line3);
nand2 M7_GSP0_SP9nc1_Xo4(M7_GSP0_SP9nc1_line2, M7_GSP0_SP9nc1_line3, M7_GSP0_line1);
inv M7_GSP0_SP9nc2_Xo0(PropXbus_4, M7_GSP0_SP9nc2_NotA);
inv M7_GSP0_SP9nc2_Xo1(M7_GSP0_line1, M7_GSP0_SP9nc2_NotB);
nand2 M7_GSP0_SP9nc2_Xo2(M7_GSP0_SP9nc2_NotA, M7_GSP0_line1, M7_GSP0_SP9nc2_line2);
nand2 M7_GSP0_SP9nc2_Xo3(M7_GSP0_SP9nc2_NotB, PropXbus_4, M7_GSP0_SP9nc2_line3);
nand2 M7_GSP0_SP9nc2_Xo4(M7_GSP0_SP9nc2_line2, M7_GSP0_SP9nc2_line3, M7_ParCin0b4_0);
inv M7_GSP1_SP9nc0_SP7c0(PropXbus_2, M7_GSP1_SP9nc0_NewInbus_6);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_0, M7_GSP1_SP9nc0_SP7c2_SP7nc0_NotA);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_1, M7_GSP1_SP9nc0_SP7c2_SP7nc0_NotB);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc0_Xo2(M7_GSP1_SP9nc0_SP7c2_SP7nc0_NotA, LocalCarryXCin1_1, M7_GSP1_SP9nc0_SP7c2_SP7nc0_line2);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc0_Xo3(M7_GSP1_SP9nc0_SP7c2_SP7nc0_NotB, LocalCarryXCin1_0, M7_GSP1_SP9nc0_SP7c2_SP7nc0_line3);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc0_Xo4(M7_GSP1_SP9nc0_SP7c2_SP7nc0_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc0_line3, M7_GSP1_SP9nc0_SP7c2_line0);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_2, M7_GSP1_SP9nc0_SP7c2_SP7nc1_NotA);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc1_Xo1(M7_GSP1_SP9nc0_SP7c2_line0, M7_GSP1_SP9nc0_SP7c2_SP7nc1_NotB);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc1_Xo2(M7_GSP1_SP9nc0_SP7c2_SP7nc1_NotA, M7_GSP1_SP9nc0_SP7c2_line0, M7_GSP1_SP9nc0_SP7c2_SP7nc1_line2);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc1_Xo3(M7_GSP1_SP9nc0_SP7c2_SP7nc1_NotB, LocalCarryXCin1_2, M7_GSP1_SP9nc0_SP7c2_SP7nc1_line3);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc1_Xo4(M7_GSP1_SP9nc0_SP7c2_SP7nc1_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc1_line3, M7_GSP1_SP9nc0_SP7c2_line1);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc2_Xo0(LocalCarryXCin1_3, M7_GSP1_SP9nc0_SP7c2_SP7nc2_NotA);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc2_Xo1(M7_GSP1_SP9nc0_SP7c2_line1, M7_GSP1_SP9nc0_SP7c2_SP7nc2_NotB);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc2_Xo2(M7_GSP1_SP9nc0_SP7c2_SP7nc2_NotA, M7_GSP1_SP9nc0_SP7c2_line1, M7_GSP1_SP9nc0_SP7c2_SP7nc2_line2);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc2_Xo3(M7_GSP1_SP9nc0_SP7c2_SP7nc2_NotB, LocalCarryXCin1_3, M7_GSP1_SP9nc0_SP7c2_SP7nc2_line3);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc2_Xo4(M7_GSP1_SP9nc0_SP7c2_SP7nc2_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc2_line3, M7_GSP1_SP9nc0_SP7c2_line2);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc3_Xo0(PropXbus_0, M7_GSP1_SP9nc0_SP7c2_SP7nc3_NotA);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc3_Xo1(M7_GSP1_SP9nc0_SP7c2_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc3_NotB);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc3_Xo2(M7_GSP1_SP9nc0_SP7c2_SP7nc3_NotA, M7_GSP1_SP9nc0_SP7c2_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc3_line2);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc3_Xo3(M7_GSP1_SP9nc0_SP7c2_SP7nc3_NotB, PropXbus_0, M7_GSP1_SP9nc0_SP7c2_SP7nc3_line3);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc3_Xo4(M7_GSP1_SP9nc0_SP7c2_SP7nc3_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc3_line3, M7_GSP1_SP9nc0_SP7c2_line3);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc4_Xo0(PropXbus_1, M7_GSP1_SP9nc0_SP7c2_SP7nc4_NotA);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc4_Xo1(M7_GSP1_SP9nc0_SP7c2_line3, M7_GSP1_SP9nc0_SP7c2_SP7nc4_NotB);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc4_Xo2(M7_GSP1_SP9nc0_SP7c2_SP7nc4_NotA, M7_GSP1_SP9nc0_SP7c2_line3, M7_GSP1_SP9nc0_SP7c2_SP7nc4_line2);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc4_Xo3(M7_GSP1_SP9nc0_SP7c2_SP7nc4_NotB, PropXbus_1, M7_GSP1_SP9nc0_SP7c2_SP7nc4_line3);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc4_Xo4(M7_GSP1_SP9nc0_SP7c2_SP7nc4_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc4_line3, M7_GSP1_SP9nc0_SP7c2_line4);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc5_Xo0(M7_GSP1_SP9nc0_NewInbus_6, M7_GSP1_SP9nc0_SP7c2_SP7nc5_NotA);
inv M7_GSP1_SP9nc0_SP7c2_SP7nc5_Xo1(M7_GSP1_SP9nc0_SP7c2_line4, M7_GSP1_SP9nc0_SP7c2_SP7nc5_NotB);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc5_Xo2(M7_GSP1_SP9nc0_SP7c2_SP7nc5_NotA, M7_GSP1_SP9nc0_SP7c2_line4, M7_GSP1_SP9nc0_SP7c2_SP7nc5_line2);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc5_Xo3(M7_GSP1_SP9nc0_SP7c2_SP7nc5_NotB, M7_GSP1_SP9nc0_NewInbus_6, M7_GSP1_SP9nc0_SP7c2_SP7nc5_line3);
nand2 M7_GSP1_SP9nc0_SP7c2_SP7nc5_Xo4(M7_GSP1_SP9nc0_SP7c2_SP7nc5_line2, M7_GSP1_SP9nc0_SP7c2_SP7nc5_line3, M7_GSP1_line0);
inv M7_GSP1_SP9nc1_Xo0(PropXbus_3, M7_GSP1_SP9nc1_NotA);
inv M7_GSP1_SP9nc1_Xo1(M7_GSP1_line0, M7_GSP1_SP9nc1_NotB);
nand2 M7_GSP1_SP9nc1_Xo2(M7_GSP1_SP9nc1_NotA, M7_GSP1_line0, M7_GSP1_SP9nc1_line2);
nand2 M7_GSP1_SP9nc1_Xo3(M7_GSP1_SP9nc1_NotB, PropXbus_3, M7_GSP1_SP9nc1_line3);
nand2 M7_GSP1_SP9nc1_Xo4(M7_GSP1_SP9nc1_line2, M7_GSP1_SP9nc1_line3, M7_GSP1_line1);
inv M7_GSP1_SP9nc2_Xo0(PropXbus_4, M7_GSP1_SP9nc2_NotA);
inv M7_GSP1_SP9nc2_Xo1(M7_GSP1_line1, M7_GSP1_SP9nc2_NotB);
nand2 M7_GSP1_SP9nc2_Xo2(M7_GSP1_SP9nc2_NotA, M7_GSP1_line1, M7_GSP1_SP9nc2_line2);
nand2 M7_GSP1_SP9nc2_Xo3(M7_GSP1_SP9nc2_NotB, PropXbus_4, M7_GSP1_SP9nc2_line3);
nand2 M7_GSP1_SP9nc2_Xo4(M7_GSP1_SP9nc2_line2, M7_GSP1_SP9nc2_line3, M7_ParCin1b4_0);
inv M7_GSP2_SP7nc0_Xo0(M5_GenXbus_5, M7_GSP2_SP7nc0_NotA);
inv M7_GSP2_SP7nc0_Xo1(LocalCarryXCin0_6, M7_GSP2_SP7nc0_NotB);
nand2 M7_GSP2_SP7nc0_Xo2(M7_GSP2_SP7nc0_NotA, LocalCarryXCin0_6, M7_GSP2_SP7nc0_line2);
nand2 M7_GSP2_SP7nc0_Xo3(M7_GSP2_SP7nc0_NotB, M5_GenXbus_5, M7_GSP2_SP7nc0_line3);
nand2 M7_GSP2_SP7nc0_Xo4(M7_GSP2_SP7nc0_line2, M7_GSP2_SP7nc0_line3, M7_GSP2_line0);
inv M7_GSP2_SP7nc1_Xo0(LocalCarryXCin0_7, M7_GSP2_SP7nc1_NotA);
inv M7_GSP2_SP7nc1_Xo1(M7_GSP2_line0, M7_GSP2_SP7nc1_NotB);
nand2 M7_GSP2_SP7nc1_Xo2(M7_GSP2_SP7nc1_NotA, M7_GSP2_line0, M7_GSP2_SP7nc1_line2);
nand2 M7_GSP2_SP7nc1_Xo3(M7_GSP2_SP7nc1_NotB, LocalCarryXCin0_7, M7_GSP2_SP7nc1_line3);
nand2 M7_GSP2_SP7nc1_Xo4(M7_GSP2_SP7nc1_line2, M7_GSP2_SP7nc1_line3, M7_GSP2_line1);
inv M7_GSP2_SP7nc2_Xo0(PropXbus_5, M7_GSP2_SP7nc2_NotA);
inv M7_GSP2_SP7nc2_Xo1(M7_GSP2_line1, M7_GSP2_SP7nc2_NotB);
nand2 M7_GSP2_SP7nc2_Xo2(M7_GSP2_SP7nc2_NotA, M7_GSP2_line1, M7_GSP2_SP7nc2_line2);
nand2 M7_GSP2_SP7nc2_Xo3(M7_GSP2_SP7nc2_NotB, PropXbus_5, M7_GSP2_SP7nc2_line3);
nand2 M7_GSP2_SP7nc2_Xo4(M7_GSP2_SP7nc2_line2, M7_GSP2_SP7nc2_line3, M7_GSP2_line2);
inv M7_GSP2_SP7nc3_Xo0(PropXbus_6, M7_GSP2_SP7nc3_NotA);
inv M7_GSP2_SP7nc3_Xo1(M7_GSP2_line2, M7_GSP2_SP7nc3_NotB);
nand2 M7_GSP2_SP7nc3_Xo2(M7_GSP2_SP7nc3_NotA, M7_GSP2_line2, M7_GSP2_SP7nc3_line2);
nand2 M7_GSP2_SP7nc3_Xo3(M7_GSP2_SP7nc3_NotB, PropXbus_6, M7_GSP2_SP7nc3_line3);
nand2 M7_GSP2_SP7nc3_Xo4(M7_GSP2_SP7nc3_line2, M7_GSP2_SP7nc3_line3, M7_GSP2_line3);
inv M7_GSP2_SP7nc4_Xo0(PropXbus_7, M7_GSP2_SP7nc4_NotA);
inv M7_GSP2_SP7nc4_Xo1(M7_GSP2_line3, M7_GSP2_SP7nc4_NotB);
nand2 M7_GSP2_SP7nc4_Xo2(M7_GSP2_SP7nc4_NotA, M7_GSP2_line3, M7_GSP2_SP7nc4_line2);
nand2 M7_GSP2_SP7nc4_Xo3(M7_GSP2_SP7nc4_NotB, PropXbus_7, M7_GSP2_SP7nc4_line3);
nand2 M7_GSP2_SP7nc4_Xo4(M7_GSP2_SP7nc4_line2, M7_GSP2_SP7nc4_line3, M7_GSP2_line4);
inv M7_GSP2_SP7nc5_Xo0(PropXbus_8, M7_GSP2_SP7nc5_NotA);
inv M7_GSP2_SP7nc5_Xo1(M7_GSP2_line4, M7_GSP2_SP7nc5_NotB);
nand2 M7_GSP2_SP7nc5_Xo2(M7_GSP2_SP7nc5_NotA, M7_GSP2_line4, M7_GSP2_SP7nc5_line2);
nand2 M7_GSP2_SP7nc5_Xo3(M7_GSP2_SP7nc5_NotB, PropXbus_8, M7_GSP2_SP7nc5_line3);
nand2 M7_GSP2_SP7nc5_Xo4(M7_GSP2_SP7nc5_line2, M7_GSP2_SP7nc5_line3, M7_ParCin0b8_5);
inv M7_GSP3_SP7c0(PropXbus_8, M7_GSP3_NewInbus_6);
inv M7_GSP3_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_5, M7_GSP3_SP7c2_SP7nc0_NotA);
inv M7_GSP3_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_6, M7_GSP3_SP7c2_SP7nc0_NotB);
nand2 M7_GSP3_SP7c2_SP7nc0_Xo2(M7_GSP3_SP7c2_SP7nc0_NotA, LocalCarryXCin1_6, M7_GSP3_SP7c2_SP7nc0_line2);
nand2 M7_GSP3_SP7c2_SP7nc0_Xo3(M7_GSP3_SP7c2_SP7nc0_NotB, LocalCarryXCin1_5, M7_GSP3_SP7c2_SP7nc0_line3);
nand2 M7_GSP3_SP7c2_SP7nc0_Xo4(M7_GSP3_SP7c2_SP7nc0_line2, M7_GSP3_SP7c2_SP7nc0_line3, M7_GSP3_SP7c2_line0);
inv M7_GSP3_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_7, M7_GSP3_SP7c2_SP7nc1_NotA);
inv M7_GSP3_SP7c2_SP7nc1_Xo1(M7_GSP3_SP7c2_line0, M7_GSP3_SP7c2_SP7nc1_NotB);
nand2 M7_GSP3_SP7c2_SP7nc1_Xo2(M7_GSP3_SP7c2_SP7nc1_NotA, M7_GSP3_SP7c2_line0, M7_GSP3_SP7c2_SP7nc1_line2);
nand2 M7_GSP3_SP7c2_SP7nc1_Xo3(M7_GSP3_SP7c2_SP7nc1_NotB, LocalCarryXCin1_7, M7_GSP3_SP7c2_SP7nc1_line3);
nand2 M7_GSP3_SP7c2_SP7nc1_Xo4(M7_GSP3_SP7c2_SP7nc1_line2, M7_GSP3_SP7c2_SP7nc1_line3, M7_GSP3_SP7c2_line1);
inv M7_GSP3_SP7c2_SP7nc2_Xo0(PropXbus_5, M7_GSP3_SP7c2_SP7nc2_NotA);
inv M7_GSP3_SP7c2_SP7nc2_Xo1(M7_GSP3_SP7c2_line1, M7_GSP3_SP7c2_SP7nc2_NotB);
nand2 M7_GSP3_SP7c2_SP7nc2_Xo2(M7_GSP3_SP7c2_SP7nc2_NotA, M7_GSP3_SP7c2_line1, M7_GSP3_SP7c2_SP7nc2_line2);
nand2 M7_GSP3_SP7c2_SP7nc2_Xo3(M7_GSP3_SP7c2_SP7nc2_NotB, PropXbus_5, M7_GSP3_SP7c2_SP7nc2_line3);
nand2 M7_GSP3_SP7c2_SP7nc2_Xo4(M7_GSP3_SP7c2_SP7nc2_line2, M7_GSP3_SP7c2_SP7nc2_line3, M7_GSP3_SP7c2_line2);
inv M7_GSP3_SP7c2_SP7nc3_Xo0(PropXbus_6, M7_GSP3_SP7c2_SP7nc3_NotA);
inv M7_GSP3_SP7c2_SP7nc3_Xo1(M7_GSP3_SP7c2_line2, M7_GSP3_SP7c2_SP7nc3_NotB);
nand2 M7_GSP3_SP7c2_SP7nc3_Xo2(M7_GSP3_SP7c2_SP7nc3_NotA, M7_GSP3_SP7c2_line2, M7_GSP3_SP7c2_SP7nc3_line2);
nand2 M7_GSP3_SP7c2_SP7nc3_Xo3(M7_GSP3_SP7c2_SP7nc3_NotB, PropXbus_6, M7_GSP3_SP7c2_SP7nc3_line3);
nand2 M7_GSP3_SP7c2_SP7nc3_Xo4(M7_GSP3_SP7c2_SP7nc3_line2, M7_GSP3_SP7c2_SP7nc3_line3, M7_GSP3_SP7c2_line3);
inv M7_GSP3_SP7c2_SP7nc4_Xo0(PropXbus_7, M7_GSP3_SP7c2_SP7nc4_NotA);
inv M7_GSP3_SP7c2_SP7nc4_Xo1(M7_GSP3_SP7c2_line3, M7_GSP3_SP7c2_SP7nc4_NotB);
nand2 M7_GSP3_SP7c2_SP7nc4_Xo2(M7_GSP3_SP7c2_SP7nc4_NotA, M7_GSP3_SP7c2_line3, M7_GSP3_SP7c2_SP7nc4_line2);
nand2 M7_GSP3_SP7c2_SP7nc4_Xo3(M7_GSP3_SP7c2_SP7nc4_NotB, PropXbus_7, M7_GSP3_SP7c2_SP7nc4_line3);
nand2 M7_GSP3_SP7c2_SP7nc4_Xo4(M7_GSP3_SP7c2_SP7nc4_line2, M7_GSP3_SP7c2_SP7nc4_line3, M7_GSP3_SP7c2_line4);
inv M7_GSP3_SP7c2_SP7nc5_Xo0(M7_GSP3_NewInbus_6, M7_GSP3_SP7c2_SP7nc5_NotA);
inv M7_GSP3_SP7c2_SP7nc5_Xo1(M7_GSP3_SP7c2_line4, M7_GSP3_SP7c2_SP7nc5_NotB);
nand2 M7_GSP3_SP7c2_SP7nc5_Xo2(M7_GSP3_SP7c2_SP7nc5_NotA, M7_GSP3_SP7c2_line4, M7_GSP3_SP7c2_SP7nc5_line2);
nand2 M7_GSP3_SP7c2_SP7nc5_Xo3(M7_GSP3_SP7c2_SP7nc5_NotB, M7_GSP3_NewInbus_6, M7_GSP3_SP7c2_SP7nc5_line3);
nand2 M7_GSP3_SP7c2_SP7nc5_Xo4(M7_GSP3_SP7c2_SP7nc5_line2, M7_GSP3_SP7c2_SP7nc5_line3, M7_ParCin1b8_5);
inv M7_GSP4_SP9nc0_SP7nc0_Xo0(M5_GenXbus_9, M7_GSP4_SP9nc0_SP7nc0_NotA);
inv M7_GSP4_SP9nc0_SP7nc0_Xo1(LocalCarryXCin0_10, M7_GSP4_SP9nc0_SP7nc0_NotB);
nand2 M7_GSP4_SP9nc0_SP7nc0_Xo2(M7_GSP4_SP9nc0_SP7nc0_NotA, LocalCarryXCin0_10, M7_GSP4_SP9nc0_SP7nc0_line2);
nand2 M7_GSP4_SP9nc0_SP7nc0_Xo3(M7_GSP4_SP9nc0_SP7nc0_NotB, M5_GenXbus_9, M7_GSP4_SP9nc0_SP7nc0_line3);
nand2 M7_GSP4_SP9nc0_SP7nc0_Xo4(M7_GSP4_SP9nc0_SP7nc0_line2, M7_GSP4_SP9nc0_SP7nc0_line3, M7_GSP4_SP9nc0_line0);
inv M7_GSP4_SP9nc0_SP7nc1_Xo0(LocalCarryXCin0_11, M7_GSP4_SP9nc0_SP7nc1_NotA);
inv M7_GSP4_SP9nc0_SP7nc1_Xo1(M7_GSP4_SP9nc0_line0, M7_GSP4_SP9nc0_SP7nc1_NotB);
nand2 M7_GSP4_SP9nc0_SP7nc1_Xo2(M7_GSP4_SP9nc0_SP7nc1_NotA, M7_GSP4_SP9nc0_line0, M7_GSP4_SP9nc0_SP7nc1_line2);
nand2 M7_GSP4_SP9nc0_SP7nc1_Xo3(M7_GSP4_SP9nc0_SP7nc1_NotB, LocalCarryXCin0_11, M7_GSP4_SP9nc0_SP7nc1_line3);
nand2 M7_GSP4_SP9nc0_SP7nc1_Xo4(M7_GSP4_SP9nc0_SP7nc1_line2, M7_GSP4_SP9nc0_SP7nc1_line3, M7_GSP4_SP9nc0_line1);
inv M7_GSP4_SP9nc0_SP7nc2_Xo0(LocalCarryXCin0_12, M7_GSP4_SP9nc0_SP7nc2_NotA);
inv M7_GSP4_SP9nc0_SP7nc2_Xo1(M7_GSP4_SP9nc0_line1, M7_GSP4_SP9nc0_SP7nc2_NotB);
nand2 M7_GSP4_SP9nc0_SP7nc2_Xo2(M7_GSP4_SP9nc0_SP7nc2_NotA, M7_GSP4_SP9nc0_line1, M7_GSP4_SP9nc0_SP7nc2_line2);
nand2 M7_GSP4_SP9nc0_SP7nc2_Xo3(M7_GSP4_SP9nc0_SP7nc2_NotB, LocalCarryXCin0_12, M7_GSP4_SP9nc0_SP7nc2_line3);
nand2 M7_GSP4_SP9nc0_SP7nc2_Xo4(M7_GSP4_SP9nc0_SP7nc2_line2, M7_GSP4_SP9nc0_SP7nc2_line3, M7_GSP4_SP9nc0_line2);
inv M7_GSP4_SP9nc0_SP7nc3_Xo0(PropXbus_9, M7_GSP4_SP9nc0_SP7nc3_NotA);
inv M7_GSP4_SP9nc0_SP7nc3_Xo1(M7_GSP4_SP9nc0_line2, M7_GSP4_SP9nc0_SP7nc3_NotB);
nand2 M7_GSP4_SP9nc0_SP7nc3_Xo2(M7_GSP4_SP9nc0_SP7nc3_NotA, M7_GSP4_SP9nc0_line2, M7_GSP4_SP9nc0_SP7nc3_line2);
nand2 M7_GSP4_SP9nc0_SP7nc3_Xo3(M7_GSP4_SP9nc0_SP7nc3_NotB, PropXbus_9, M7_GSP4_SP9nc0_SP7nc3_line3);
nand2 M7_GSP4_SP9nc0_SP7nc3_Xo4(M7_GSP4_SP9nc0_SP7nc3_line2, M7_GSP4_SP9nc0_SP7nc3_line3, M7_GSP4_SP9nc0_line3);
inv M7_GSP4_SP9nc0_SP7nc4_Xo0(PropXbus_10, M7_GSP4_SP9nc0_SP7nc4_NotA);
inv M7_GSP4_SP9nc0_SP7nc4_Xo1(M7_GSP4_SP9nc0_line3, M7_GSP4_SP9nc0_SP7nc4_NotB);
nand2 M7_GSP4_SP9nc0_SP7nc4_Xo2(M7_GSP4_SP9nc0_SP7nc4_NotA, M7_GSP4_SP9nc0_line3, M7_GSP4_SP9nc0_SP7nc4_line2);
nand2 M7_GSP4_SP9nc0_SP7nc4_Xo3(M7_GSP4_SP9nc0_SP7nc4_NotB, PropXbus_10, M7_GSP4_SP9nc0_SP7nc4_line3);
nand2 M7_GSP4_SP9nc0_SP7nc4_Xo4(M7_GSP4_SP9nc0_SP7nc4_line2, M7_GSP4_SP9nc0_SP7nc4_line3, M7_GSP4_SP9nc0_line4);
inv M7_GSP4_SP9nc0_SP7nc5_Xo0(PropXbus_11, M7_GSP4_SP9nc0_SP7nc5_NotA);
inv M7_GSP4_SP9nc0_SP7nc5_Xo1(M7_GSP4_SP9nc0_line4, M7_GSP4_SP9nc0_SP7nc5_NotB);
nand2 M7_GSP4_SP9nc0_SP7nc5_Xo2(M7_GSP4_SP9nc0_SP7nc5_NotA, M7_GSP4_SP9nc0_line4, M7_GSP4_SP9nc0_SP7nc5_line2);
nand2 M7_GSP4_SP9nc0_SP7nc5_Xo3(M7_GSP4_SP9nc0_SP7nc5_NotB, PropXbus_11, M7_GSP4_SP9nc0_SP7nc5_line3);
nand2 M7_GSP4_SP9nc0_SP7nc5_Xo4(M7_GSP4_SP9nc0_SP7nc5_line2, M7_GSP4_SP9nc0_SP7nc5_line3, M7_GSP4_line0);
inv M7_GSP4_SP9nc1_Xo0(PropXbus_12, M7_GSP4_SP9nc1_NotA);
inv M7_GSP4_SP9nc1_Xo1(M7_GSP4_line0, M7_GSP4_SP9nc1_NotB);
nand2 M7_GSP4_SP9nc1_Xo2(M7_GSP4_SP9nc1_NotA, M7_GSP4_line0, M7_GSP4_SP9nc1_line2);
nand2 M7_GSP4_SP9nc1_Xo3(M7_GSP4_SP9nc1_NotB, PropXbus_12, M7_GSP4_SP9nc1_line3);
nand2 M7_GSP4_SP9nc1_Xo4(M7_GSP4_SP9nc1_line2, M7_GSP4_SP9nc1_line3, M7_GSP4_line1);
inv M7_GSP4_SP9nc2_Xo0(PropXbus_13, M7_GSP4_SP9nc2_NotA);
inv M7_GSP4_SP9nc2_Xo1(M7_GSP4_line1, M7_GSP4_SP9nc2_NotB);
nand2 M7_GSP4_SP9nc2_Xo2(M7_GSP4_SP9nc2_NotA, M7_GSP4_line1, M7_GSP4_SP9nc2_line2);
nand2 M7_GSP4_SP9nc2_Xo3(M7_GSP4_SP9nc2_NotB, PropXbus_13, M7_GSP4_SP9nc2_line3);
nand2 M7_GSP4_SP9nc2_Xo4(M7_GSP4_SP9nc2_line2, M7_GSP4_SP9nc2_line3, M7_ParCin0b13_9);
inv M7_GSP5_SP9nc0_SP7c0(PropXbus_11, M7_GSP5_SP9nc0_NewInbus_6);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_9, M7_GSP5_SP9nc0_SP7c2_SP7nc0_NotA);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_10, M7_GSP5_SP9nc0_SP7c2_SP7nc0_NotB);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc0_Xo2(M7_GSP5_SP9nc0_SP7c2_SP7nc0_NotA, LocalCarryXCin1_10, M7_GSP5_SP9nc0_SP7c2_SP7nc0_line2);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc0_Xo3(M7_GSP5_SP9nc0_SP7c2_SP7nc0_NotB, LocalCarryXCin1_9, M7_GSP5_SP9nc0_SP7c2_SP7nc0_line3);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc0_Xo4(M7_GSP5_SP9nc0_SP7c2_SP7nc0_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc0_line3, M7_GSP5_SP9nc0_SP7c2_line0);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_11, M7_GSP5_SP9nc0_SP7c2_SP7nc1_NotA);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc1_Xo1(M7_GSP5_SP9nc0_SP7c2_line0, M7_GSP5_SP9nc0_SP7c2_SP7nc1_NotB);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc1_Xo2(M7_GSP5_SP9nc0_SP7c2_SP7nc1_NotA, M7_GSP5_SP9nc0_SP7c2_line0, M7_GSP5_SP9nc0_SP7c2_SP7nc1_line2);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc1_Xo3(M7_GSP5_SP9nc0_SP7c2_SP7nc1_NotB, LocalCarryXCin1_11, M7_GSP5_SP9nc0_SP7c2_SP7nc1_line3);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc1_Xo4(M7_GSP5_SP9nc0_SP7c2_SP7nc1_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc1_line3, M7_GSP5_SP9nc0_SP7c2_line1);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc2_Xo0(LocalCarryXCin1_12, M7_GSP5_SP9nc0_SP7c2_SP7nc2_NotA);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc2_Xo1(M7_GSP5_SP9nc0_SP7c2_line1, M7_GSP5_SP9nc0_SP7c2_SP7nc2_NotB);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc2_Xo2(M7_GSP5_SP9nc0_SP7c2_SP7nc2_NotA, M7_GSP5_SP9nc0_SP7c2_line1, M7_GSP5_SP9nc0_SP7c2_SP7nc2_line2);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc2_Xo3(M7_GSP5_SP9nc0_SP7c2_SP7nc2_NotB, LocalCarryXCin1_12, M7_GSP5_SP9nc0_SP7c2_SP7nc2_line3);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc2_Xo4(M7_GSP5_SP9nc0_SP7c2_SP7nc2_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc2_line3, M7_GSP5_SP9nc0_SP7c2_line2);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc3_Xo0(PropXbus_9, M7_GSP5_SP9nc0_SP7c2_SP7nc3_NotA);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc3_Xo1(M7_GSP5_SP9nc0_SP7c2_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc3_NotB);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc3_Xo2(M7_GSP5_SP9nc0_SP7c2_SP7nc3_NotA, M7_GSP5_SP9nc0_SP7c2_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc3_line2);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc3_Xo3(M7_GSP5_SP9nc0_SP7c2_SP7nc3_NotB, PropXbus_9, M7_GSP5_SP9nc0_SP7c2_SP7nc3_line3);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc3_Xo4(M7_GSP5_SP9nc0_SP7c2_SP7nc3_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc3_line3, M7_GSP5_SP9nc0_SP7c2_line3);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc4_Xo0(PropXbus_10, M7_GSP5_SP9nc0_SP7c2_SP7nc4_NotA);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc4_Xo1(M7_GSP5_SP9nc0_SP7c2_line3, M7_GSP5_SP9nc0_SP7c2_SP7nc4_NotB);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc4_Xo2(M7_GSP5_SP9nc0_SP7c2_SP7nc4_NotA, M7_GSP5_SP9nc0_SP7c2_line3, M7_GSP5_SP9nc0_SP7c2_SP7nc4_line2);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc4_Xo3(M7_GSP5_SP9nc0_SP7c2_SP7nc4_NotB, PropXbus_10, M7_GSP5_SP9nc0_SP7c2_SP7nc4_line3);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc4_Xo4(M7_GSP5_SP9nc0_SP7c2_SP7nc4_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc4_line3, M7_GSP5_SP9nc0_SP7c2_line4);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc5_Xo0(M7_GSP5_SP9nc0_NewInbus_6, M7_GSP5_SP9nc0_SP7c2_SP7nc5_NotA);
inv M7_GSP5_SP9nc0_SP7c2_SP7nc5_Xo1(M7_GSP5_SP9nc0_SP7c2_line4, M7_GSP5_SP9nc0_SP7c2_SP7nc5_NotB);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc5_Xo2(M7_GSP5_SP9nc0_SP7c2_SP7nc5_NotA, M7_GSP5_SP9nc0_SP7c2_line4, M7_GSP5_SP9nc0_SP7c2_SP7nc5_line2);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc5_Xo3(M7_GSP5_SP9nc0_SP7c2_SP7nc5_NotB, M7_GSP5_SP9nc0_NewInbus_6, M7_GSP5_SP9nc0_SP7c2_SP7nc5_line3);
nand2 M7_GSP5_SP9nc0_SP7c2_SP7nc5_Xo4(M7_GSP5_SP9nc0_SP7c2_SP7nc5_line2, M7_GSP5_SP9nc0_SP7c2_SP7nc5_line3, M7_GSP5_line0);
inv M7_GSP5_SP9nc1_Xo0(PropXbus_12, M7_GSP5_SP9nc1_NotA);
inv M7_GSP5_SP9nc1_Xo1(M7_GSP5_line0, M7_GSP5_SP9nc1_NotB);
nand2 M7_GSP5_SP9nc1_Xo2(M7_GSP5_SP9nc1_NotA, M7_GSP5_line0, M7_GSP5_SP9nc1_line2);
nand2 M7_GSP5_SP9nc1_Xo3(M7_GSP5_SP9nc1_NotB, PropXbus_12, M7_GSP5_SP9nc1_line3);
nand2 M7_GSP5_SP9nc1_Xo4(M7_GSP5_SP9nc1_line2, M7_GSP5_SP9nc1_line3, M7_GSP5_line1);
inv M7_GSP5_SP9nc2_Xo0(PropXbus_13, M7_GSP5_SP9nc2_NotA);
inv M7_GSP5_SP9nc2_Xo1(M7_GSP5_line1, M7_GSP5_SP9nc2_NotB);
nand2 M7_GSP5_SP9nc2_Xo2(M7_GSP5_SP9nc2_NotA, M7_GSP5_line1, M7_GSP5_SP9nc2_line2);
nand2 M7_GSP5_SP9nc2_Xo3(M7_GSP5_SP9nc2_NotB, PropXbus_13, M7_GSP5_SP9nc2_line3);
nand2 M7_GSP5_SP9nc2_Xo4(M7_GSP5_SP9nc2_line2, M7_GSP5_SP9nc2_line3, M7_ParCin1b13_9);
inv M7_GSP6_SP7nc0_Xo0(M5_GenXbus_14, M7_GSP6_SP7nc0_NotA);
inv M7_GSP6_SP7nc0_Xo1(LocalCarryXCin0_15, M7_GSP6_SP7nc0_NotB);
nand2 M7_GSP6_SP7nc0_Xo2(M7_GSP6_SP7nc0_NotA, LocalCarryXCin0_15, M7_GSP6_SP7nc0_line2);
nand2 M7_GSP6_SP7nc0_Xo3(M7_GSP6_SP7nc0_NotB, M5_GenXbus_14, M7_GSP6_SP7nc0_line3);
nand2 M7_GSP6_SP7nc0_Xo4(M7_GSP6_SP7nc0_line2, M7_GSP6_SP7nc0_line3, M7_GSP6_line0);
inv M7_GSP6_SP7nc1_Xo0(LocalCarryXCin0_16, M7_GSP6_SP7nc1_NotA);
inv M7_GSP6_SP7nc1_Xo1(M7_GSP6_line0, M7_GSP6_SP7nc1_NotB);
nand2 M7_GSP6_SP7nc1_Xo2(M7_GSP6_SP7nc1_NotA, M7_GSP6_line0, M7_GSP6_SP7nc1_line2);
nand2 M7_GSP6_SP7nc1_Xo3(M7_GSP6_SP7nc1_NotB, LocalCarryXCin0_16, M7_GSP6_SP7nc1_line3);
nand2 M7_GSP6_SP7nc1_Xo4(M7_GSP6_SP7nc1_line2, M7_GSP6_SP7nc1_line3, M7_GSP6_line1);
inv M7_GSP6_SP7nc2_Xo0(PropXbus_14, M7_GSP6_SP7nc2_NotA);
inv M7_GSP6_SP7nc2_Xo1(M7_GSP6_line1, M7_GSP6_SP7nc2_NotB);
nand2 M7_GSP6_SP7nc2_Xo2(M7_GSP6_SP7nc2_NotA, M7_GSP6_line1, M7_GSP6_SP7nc2_line2);
nand2 M7_GSP6_SP7nc2_Xo3(M7_GSP6_SP7nc2_NotB, PropXbus_14, M7_GSP6_SP7nc2_line3);
nand2 M7_GSP6_SP7nc2_Xo4(M7_GSP6_SP7nc2_line2, M7_GSP6_SP7nc2_line3, M7_GSP6_line2);
inv M7_GSP6_SP7nc3_Xo0(PropXbus_15, M7_GSP6_SP7nc3_NotA);
inv M7_GSP6_SP7nc3_Xo1(M7_GSP6_line2, M7_GSP6_SP7nc3_NotB);
nand2 M7_GSP6_SP7nc3_Xo2(M7_GSP6_SP7nc3_NotA, M7_GSP6_line2, M7_GSP6_SP7nc3_line2);
nand2 M7_GSP6_SP7nc3_Xo3(M7_GSP6_SP7nc3_NotB, PropXbus_15, M7_GSP6_SP7nc3_line3);
nand2 M7_GSP6_SP7nc3_Xo4(M7_GSP6_SP7nc3_line2, M7_GSP6_SP7nc3_line3, M7_GSP6_line3);
inv M7_GSP6_SP7nc4_Xo0(PropXbus_16, M7_GSP6_SP7nc4_NotA);
inv M7_GSP6_SP7nc4_Xo1(M7_GSP6_line3, M7_GSP6_SP7nc4_NotB);
nand2 M7_GSP6_SP7nc4_Xo2(M7_GSP6_SP7nc4_NotA, M7_GSP6_line3, M7_GSP6_SP7nc4_line2);
nand2 M7_GSP6_SP7nc4_Xo3(M7_GSP6_SP7nc4_NotB, PropXbus_16, M7_GSP6_SP7nc4_line3);
nand2 M7_GSP6_SP7nc4_Xo4(M7_GSP6_SP7nc4_line2, M7_GSP6_SP7nc4_line3, M7_GSP6_line4);
inv M7_GSP6_SP7nc5_Xo0(PropXbus_17, M7_GSP6_SP7nc5_NotA);
inv M7_GSP6_SP7nc5_Xo1(M7_GSP6_line4, M7_GSP6_SP7nc5_NotB);
nand2 M7_GSP6_SP7nc5_Xo2(M7_GSP6_SP7nc5_NotA, M7_GSP6_line4, M7_GSP6_SP7nc5_line2);
nand2 M7_GSP6_SP7nc5_Xo3(M7_GSP6_SP7nc5_NotB, PropXbus_17, M7_GSP6_SP7nc5_line3);
nand2 M7_GSP6_SP7nc5_Xo4(M7_GSP6_SP7nc5_line2, M7_GSP6_SP7nc5_line3, M7_ParCin0b17_14);
inv M7_GSP7_SP7c0(PropXbus_17, M7_GSP7_NewInbus_6);
inv M7_GSP7_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_14, M7_GSP7_SP7c2_SP7nc0_NotA);
inv M7_GSP7_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_15, M7_GSP7_SP7c2_SP7nc0_NotB);
nand2 M7_GSP7_SP7c2_SP7nc0_Xo2(M7_GSP7_SP7c2_SP7nc0_NotA, LocalCarryXCin1_15, M7_GSP7_SP7c2_SP7nc0_line2);
nand2 M7_GSP7_SP7c2_SP7nc0_Xo3(M7_GSP7_SP7c2_SP7nc0_NotB, LocalCarryXCin1_14, M7_GSP7_SP7c2_SP7nc0_line3);
nand2 M7_GSP7_SP7c2_SP7nc0_Xo4(M7_GSP7_SP7c2_SP7nc0_line2, M7_GSP7_SP7c2_SP7nc0_line3, M7_GSP7_SP7c2_line0);
inv M7_GSP7_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_16, M7_GSP7_SP7c2_SP7nc1_NotA);
inv M7_GSP7_SP7c2_SP7nc1_Xo1(M7_GSP7_SP7c2_line0, M7_GSP7_SP7c2_SP7nc1_NotB);
nand2 M7_GSP7_SP7c2_SP7nc1_Xo2(M7_GSP7_SP7c2_SP7nc1_NotA, M7_GSP7_SP7c2_line0, M7_GSP7_SP7c2_SP7nc1_line2);
nand2 M7_GSP7_SP7c2_SP7nc1_Xo3(M7_GSP7_SP7c2_SP7nc1_NotB, LocalCarryXCin1_16, M7_GSP7_SP7c2_SP7nc1_line3);
nand2 M7_GSP7_SP7c2_SP7nc1_Xo4(M7_GSP7_SP7c2_SP7nc1_line2, M7_GSP7_SP7c2_SP7nc1_line3, M7_GSP7_SP7c2_line1);
inv M7_GSP7_SP7c2_SP7nc2_Xo0(PropXbus_14, M7_GSP7_SP7c2_SP7nc2_NotA);
inv M7_GSP7_SP7c2_SP7nc2_Xo1(M7_GSP7_SP7c2_line1, M7_GSP7_SP7c2_SP7nc2_NotB);
nand2 M7_GSP7_SP7c2_SP7nc2_Xo2(M7_GSP7_SP7c2_SP7nc2_NotA, M7_GSP7_SP7c2_line1, M7_GSP7_SP7c2_SP7nc2_line2);
nand2 M7_GSP7_SP7c2_SP7nc2_Xo3(M7_GSP7_SP7c2_SP7nc2_NotB, PropXbus_14, M7_GSP7_SP7c2_SP7nc2_line3);
nand2 M7_GSP7_SP7c2_SP7nc2_Xo4(M7_GSP7_SP7c2_SP7nc2_line2, M7_GSP7_SP7c2_SP7nc2_line3, M7_GSP7_SP7c2_line2);
inv M7_GSP7_SP7c2_SP7nc3_Xo0(PropXbus_15, M7_GSP7_SP7c2_SP7nc3_NotA);
inv M7_GSP7_SP7c2_SP7nc3_Xo1(M7_GSP7_SP7c2_line2, M7_GSP7_SP7c2_SP7nc3_NotB);
nand2 M7_GSP7_SP7c2_SP7nc3_Xo2(M7_GSP7_SP7c2_SP7nc3_NotA, M7_GSP7_SP7c2_line2, M7_GSP7_SP7c2_SP7nc3_line2);
nand2 M7_GSP7_SP7c2_SP7nc3_Xo3(M7_GSP7_SP7c2_SP7nc3_NotB, PropXbus_15, M7_GSP7_SP7c2_SP7nc3_line3);
nand2 M7_GSP7_SP7c2_SP7nc3_Xo4(M7_GSP7_SP7c2_SP7nc3_line2, M7_GSP7_SP7c2_SP7nc3_line3, M7_GSP7_SP7c2_line3);
inv M7_GSP7_SP7c2_SP7nc4_Xo0(PropXbus_16, M7_GSP7_SP7c2_SP7nc4_NotA);
inv M7_GSP7_SP7c2_SP7nc4_Xo1(M7_GSP7_SP7c2_line3, M7_GSP7_SP7c2_SP7nc4_NotB);
nand2 M7_GSP7_SP7c2_SP7nc4_Xo2(M7_GSP7_SP7c2_SP7nc4_NotA, M7_GSP7_SP7c2_line3, M7_GSP7_SP7c2_SP7nc4_line2);
nand2 M7_GSP7_SP7c2_SP7nc4_Xo3(M7_GSP7_SP7c2_SP7nc4_NotB, PropXbus_16, M7_GSP7_SP7c2_SP7nc4_line3);
nand2 M7_GSP7_SP7c2_SP7nc4_Xo4(M7_GSP7_SP7c2_SP7nc4_line2, M7_GSP7_SP7c2_SP7nc4_line3, M7_GSP7_SP7c2_line4);
inv M7_GSP7_SP7c2_SP7nc5_Xo0(M7_GSP7_NewInbus_6, M7_GSP7_SP7c2_SP7nc5_NotA);
inv M7_GSP7_SP7c2_SP7nc5_Xo1(M7_GSP7_SP7c2_line4, M7_GSP7_SP7c2_SP7nc5_NotB);
nand2 M7_GSP7_SP7c2_SP7nc5_Xo2(M7_GSP7_SP7c2_SP7nc5_NotA, M7_GSP7_SP7c2_line4, M7_GSP7_SP7c2_SP7nc5_line2);
nand2 M7_GSP7_SP7c2_SP7nc5_Xo3(M7_GSP7_SP7c2_SP7nc5_NotB, M7_GSP7_NewInbus_6, M7_GSP7_SP7c2_SP7nc5_line3);
nand2 M7_GSP7_SP7c2_SP7nc5_Xo4(M7_GSP7_SP7c2_SP7nc5_line2, M7_GSP7_SP7c2_SP7nc5_line3, M7_ParCin1b17_14);
inv M7_GSP8_SP9nc0_SP7nc0_Xo0(M5_GenXbus_18, M7_GSP8_SP9nc0_SP7nc0_NotA);
inv M7_GSP8_SP9nc0_SP7nc0_Xo1(LocalCarryXCin0_19, M7_GSP8_SP9nc0_SP7nc0_NotB);
nand2 M7_GSP8_SP9nc0_SP7nc0_Xo2(M7_GSP8_SP9nc0_SP7nc0_NotA, LocalCarryXCin0_19, M7_GSP8_SP9nc0_SP7nc0_line2);
nand2 M7_GSP8_SP9nc0_SP7nc0_Xo3(M7_GSP8_SP9nc0_SP7nc0_NotB, M5_GenXbus_18, M7_GSP8_SP9nc0_SP7nc0_line3);
nand2 M7_GSP8_SP9nc0_SP7nc0_Xo4(M7_GSP8_SP9nc0_SP7nc0_line2, M7_GSP8_SP9nc0_SP7nc0_line3, M7_GSP8_SP9nc0_line0);
inv M7_GSP8_SP9nc0_SP7nc1_Xo0(LocalCarryXCin0_20, M7_GSP8_SP9nc0_SP7nc1_NotA);
inv M7_GSP8_SP9nc0_SP7nc1_Xo1(M7_GSP8_SP9nc0_line0, M7_GSP8_SP9nc0_SP7nc1_NotB);
nand2 M7_GSP8_SP9nc0_SP7nc1_Xo2(M7_GSP8_SP9nc0_SP7nc1_NotA, M7_GSP8_SP9nc0_line0, M7_GSP8_SP9nc0_SP7nc1_line2);
nand2 M7_GSP8_SP9nc0_SP7nc1_Xo3(M7_GSP8_SP9nc0_SP7nc1_NotB, LocalCarryXCin0_20, M7_GSP8_SP9nc0_SP7nc1_line3);
nand2 M7_GSP8_SP9nc0_SP7nc1_Xo4(M7_GSP8_SP9nc0_SP7nc1_line2, M7_GSP8_SP9nc0_SP7nc1_line3, M7_GSP8_SP9nc0_line1);
inv M7_GSP8_SP9nc0_SP7nc2_Xo0(LocalCarryXCin0_21, M7_GSP8_SP9nc0_SP7nc2_NotA);
inv M7_GSP8_SP9nc0_SP7nc2_Xo1(M7_GSP8_SP9nc0_line1, M7_GSP8_SP9nc0_SP7nc2_NotB);
nand2 M7_GSP8_SP9nc0_SP7nc2_Xo2(M7_GSP8_SP9nc0_SP7nc2_NotA, M7_GSP8_SP9nc0_line1, M7_GSP8_SP9nc0_SP7nc2_line2);
nand2 M7_GSP8_SP9nc0_SP7nc2_Xo3(M7_GSP8_SP9nc0_SP7nc2_NotB, LocalCarryXCin0_21, M7_GSP8_SP9nc0_SP7nc2_line3);
nand2 M7_GSP8_SP9nc0_SP7nc2_Xo4(M7_GSP8_SP9nc0_SP7nc2_line2, M7_GSP8_SP9nc0_SP7nc2_line3, M7_GSP8_SP9nc0_line2);
inv M7_GSP8_SP9nc0_SP7nc3_Xo0(PropXbus_18, M7_GSP8_SP9nc0_SP7nc3_NotA);
inv M7_GSP8_SP9nc0_SP7nc3_Xo1(M7_GSP8_SP9nc0_line2, M7_GSP8_SP9nc0_SP7nc3_NotB);
nand2 M7_GSP8_SP9nc0_SP7nc3_Xo2(M7_GSP8_SP9nc0_SP7nc3_NotA, M7_GSP8_SP9nc0_line2, M7_GSP8_SP9nc0_SP7nc3_line2);
nand2 M7_GSP8_SP9nc0_SP7nc3_Xo3(M7_GSP8_SP9nc0_SP7nc3_NotB, PropXbus_18, M7_GSP8_SP9nc0_SP7nc3_line3);
nand2 M7_GSP8_SP9nc0_SP7nc3_Xo4(M7_GSP8_SP9nc0_SP7nc3_line2, M7_GSP8_SP9nc0_SP7nc3_line3, M7_GSP8_SP9nc0_line3);
inv M7_GSP8_SP9nc0_SP7nc4_Xo0(PropXbus_19, M7_GSP8_SP9nc0_SP7nc4_NotA);
inv M7_GSP8_SP9nc0_SP7nc4_Xo1(M7_GSP8_SP9nc0_line3, M7_GSP8_SP9nc0_SP7nc4_NotB);
nand2 M7_GSP8_SP9nc0_SP7nc4_Xo2(M7_GSP8_SP9nc0_SP7nc4_NotA, M7_GSP8_SP9nc0_line3, M7_GSP8_SP9nc0_SP7nc4_line2);
nand2 M7_GSP8_SP9nc0_SP7nc4_Xo3(M7_GSP8_SP9nc0_SP7nc4_NotB, PropXbus_19, M7_GSP8_SP9nc0_SP7nc4_line3);
nand2 M7_GSP8_SP9nc0_SP7nc4_Xo4(M7_GSP8_SP9nc0_SP7nc4_line2, M7_GSP8_SP9nc0_SP7nc4_line3, M7_GSP8_SP9nc0_line4);
inv M7_GSP8_SP9nc0_SP7nc5_Xo0(PropXbus_20, M7_GSP8_SP9nc0_SP7nc5_NotA);
inv M7_GSP8_SP9nc0_SP7nc5_Xo1(M7_GSP8_SP9nc0_line4, M7_GSP8_SP9nc0_SP7nc5_NotB);
nand2 M7_GSP8_SP9nc0_SP7nc5_Xo2(M7_GSP8_SP9nc0_SP7nc5_NotA, M7_GSP8_SP9nc0_line4, M7_GSP8_SP9nc0_SP7nc5_line2);
nand2 M7_GSP8_SP9nc0_SP7nc5_Xo3(M7_GSP8_SP9nc0_SP7nc5_NotB, PropXbus_20, M7_GSP8_SP9nc0_SP7nc5_line3);
nand2 M7_GSP8_SP9nc0_SP7nc5_Xo4(M7_GSP8_SP9nc0_SP7nc5_line2, M7_GSP8_SP9nc0_SP7nc5_line3, M7_GSP8_line0);
inv M7_GSP8_SP9nc1_Xo0(PropXbus_21, M7_GSP8_SP9nc1_NotA);
inv M7_GSP8_SP9nc1_Xo1(M7_GSP8_line0, M7_GSP8_SP9nc1_NotB);
nand2 M7_GSP8_SP9nc1_Xo2(M7_GSP8_SP9nc1_NotA, M7_GSP8_line0, M7_GSP8_SP9nc1_line2);
nand2 M7_GSP8_SP9nc1_Xo3(M7_GSP8_SP9nc1_NotB, PropXbus_21, M7_GSP8_SP9nc1_line3);
nand2 M7_GSP8_SP9nc1_Xo4(M7_GSP8_SP9nc1_line2, M7_GSP8_SP9nc1_line3, M7_GSP8_line1);
inv M7_GSP8_SP9nc2_Xo0(PropXbus_22, M7_GSP8_SP9nc2_NotA);
inv M7_GSP8_SP9nc2_Xo1(M7_GSP8_line1, M7_GSP8_SP9nc2_NotB);
nand2 M7_GSP8_SP9nc2_Xo2(M7_GSP8_SP9nc2_NotA, M7_GSP8_line1, M7_GSP8_SP9nc2_line2);
nand2 M7_GSP8_SP9nc2_Xo3(M7_GSP8_SP9nc2_NotB, PropXbus_22, M7_GSP8_SP9nc2_line3);
nand2 M7_GSP8_SP9nc2_Xo4(M7_GSP8_SP9nc2_line2, M7_GSP8_SP9nc2_line3, M7_ParCin0b22_18);
inv M7_GSP9_SP9nc0_SP7c0(PropXbus_20, M7_GSP9_SP9nc0_NewInbus_6);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_18, M7_GSP9_SP9nc0_SP7c2_SP7nc0_NotA);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_19, M7_GSP9_SP9nc0_SP7c2_SP7nc0_NotB);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc0_Xo2(M7_GSP9_SP9nc0_SP7c2_SP7nc0_NotA, LocalCarryXCin1_19, M7_GSP9_SP9nc0_SP7c2_SP7nc0_line2);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc0_Xo3(M7_GSP9_SP9nc0_SP7c2_SP7nc0_NotB, LocalCarryXCin1_18, M7_GSP9_SP9nc0_SP7c2_SP7nc0_line3);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc0_Xo4(M7_GSP9_SP9nc0_SP7c2_SP7nc0_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc0_line3, M7_GSP9_SP9nc0_SP7c2_line0);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_20, M7_GSP9_SP9nc0_SP7c2_SP7nc1_NotA);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc1_Xo1(M7_GSP9_SP9nc0_SP7c2_line0, M7_GSP9_SP9nc0_SP7c2_SP7nc1_NotB);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc1_Xo2(M7_GSP9_SP9nc0_SP7c2_SP7nc1_NotA, M7_GSP9_SP9nc0_SP7c2_line0, M7_GSP9_SP9nc0_SP7c2_SP7nc1_line2);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc1_Xo3(M7_GSP9_SP9nc0_SP7c2_SP7nc1_NotB, LocalCarryXCin1_20, M7_GSP9_SP9nc0_SP7c2_SP7nc1_line3);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc1_Xo4(M7_GSP9_SP9nc0_SP7c2_SP7nc1_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc1_line3, M7_GSP9_SP9nc0_SP7c2_line1);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc2_Xo0(LocalCarryXCin1_21, M7_GSP9_SP9nc0_SP7c2_SP7nc2_NotA);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc2_Xo1(M7_GSP9_SP9nc0_SP7c2_line1, M7_GSP9_SP9nc0_SP7c2_SP7nc2_NotB);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc2_Xo2(M7_GSP9_SP9nc0_SP7c2_SP7nc2_NotA, M7_GSP9_SP9nc0_SP7c2_line1, M7_GSP9_SP9nc0_SP7c2_SP7nc2_line2);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc2_Xo3(M7_GSP9_SP9nc0_SP7c2_SP7nc2_NotB, LocalCarryXCin1_21, M7_GSP9_SP9nc0_SP7c2_SP7nc2_line3);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc2_Xo4(M7_GSP9_SP9nc0_SP7c2_SP7nc2_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc2_line3, M7_GSP9_SP9nc0_SP7c2_line2);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc3_Xo0(PropXbus_18, M7_GSP9_SP9nc0_SP7c2_SP7nc3_NotA);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc3_Xo1(M7_GSP9_SP9nc0_SP7c2_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc3_NotB);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc3_Xo2(M7_GSP9_SP9nc0_SP7c2_SP7nc3_NotA, M7_GSP9_SP9nc0_SP7c2_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc3_line2);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc3_Xo3(M7_GSP9_SP9nc0_SP7c2_SP7nc3_NotB, PropXbus_18, M7_GSP9_SP9nc0_SP7c2_SP7nc3_line3);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc3_Xo4(M7_GSP9_SP9nc0_SP7c2_SP7nc3_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc3_line3, M7_GSP9_SP9nc0_SP7c2_line3);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc4_Xo0(PropXbus_19, M7_GSP9_SP9nc0_SP7c2_SP7nc4_NotA);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc4_Xo1(M7_GSP9_SP9nc0_SP7c2_line3, M7_GSP9_SP9nc0_SP7c2_SP7nc4_NotB);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc4_Xo2(M7_GSP9_SP9nc0_SP7c2_SP7nc4_NotA, M7_GSP9_SP9nc0_SP7c2_line3, M7_GSP9_SP9nc0_SP7c2_SP7nc4_line2);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc4_Xo3(M7_GSP9_SP9nc0_SP7c2_SP7nc4_NotB, PropXbus_19, M7_GSP9_SP9nc0_SP7c2_SP7nc4_line3);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc4_Xo4(M7_GSP9_SP9nc0_SP7c2_SP7nc4_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc4_line3, M7_GSP9_SP9nc0_SP7c2_line4);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc5_Xo0(M7_GSP9_SP9nc0_NewInbus_6, M7_GSP9_SP9nc0_SP7c2_SP7nc5_NotA);
inv M7_GSP9_SP9nc0_SP7c2_SP7nc5_Xo1(M7_GSP9_SP9nc0_SP7c2_line4, M7_GSP9_SP9nc0_SP7c2_SP7nc5_NotB);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc5_Xo2(M7_GSP9_SP9nc0_SP7c2_SP7nc5_NotA, M7_GSP9_SP9nc0_SP7c2_line4, M7_GSP9_SP9nc0_SP7c2_SP7nc5_line2);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc5_Xo3(M7_GSP9_SP9nc0_SP7c2_SP7nc5_NotB, M7_GSP9_SP9nc0_NewInbus_6, M7_GSP9_SP9nc0_SP7c2_SP7nc5_line3);
nand2 M7_GSP9_SP9nc0_SP7c2_SP7nc5_Xo4(M7_GSP9_SP9nc0_SP7c2_SP7nc5_line2, M7_GSP9_SP9nc0_SP7c2_SP7nc5_line3, M7_GSP9_line0);
inv M7_GSP9_SP9nc1_Xo0(PropXbus_21, M7_GSP9_SP9nc1_NotA);
inv M7_GSP9_SP9nc1_Xo1(M7_GSP9_line0, M7_GSP9_SP9nc1_NotB);
nand2 M7_GSP9_SP9nc1_Xo2(M7_GSP9_SP9nc1_NotA, M7_GSP9_line0, M7_GSP9_SP9nc1_line2);
nand2 M7_GSP9_SP9nc1_Xo3(M7_GSP9_SP9nc1_NotB, PropXbus_21, M7_GSP9_SP9nc1_line3);
nand2 M7_GSP9_SP9nc1_Xo4(M7_GSP9_SP9nc1_line2, M7_GSP9_SP9nc1_line3, M7_GSP9_line1);
inv M7_GSP9_SP9nc2_Xo0(PropXbus_22, M7_GSP9_SP9nc2_NotA);
inv M7_GSP9_SP9nc2_Xo1(M7_GSP9_line1, M7_GSP9_SP9nc2_NotB);
nand2 M7_GSP9_SP9nc2_Xo2(M7_GSP9_SP9nc2_NotA, M7_GSP9_line1, M7_GSP9_SP9nc2_line2);
nand2 M7_GSP9_SP9nc2_Xo3(M7_GSP9_SP9nc2_NotB, PropXbus_22, M7_GSP9_SP9nc2_line3);
nand2 M7_GSP9_SP9nc2_Xo4(M7_GSP9_SP9nc2_line2, M7_GSP9_SP9nc2_line3, M7_ParCin1b22_18);
inv M7_GSP10_SP7nc0_Xo0(M5_GenXbus_23, M7_GSP10_SP7nc0_NotA);
inv M7_GSP10_SP7nc0_Xo1(LocalCarryXCin0_24, M7_GSP10_SP7nc0_NotB);
nand2 M7_GSP10_SP7nc0_Xo2(M7_GSP10_SP7nc0_NotA, LocalCarryXCin0_24, M7_GSP10_SP7nc0_line2);
nand2 M7_GSP10_SP7nc0_Xo3(M7_GSP10_SP7nc0_NotB, M5_GenXbus_23, M7_GSP10_SP7nc0_line3);
nand2 M7_GSP10_SP7nc0_Xo4(M7_GSP10_SP7nc0_line2, M7_GSP10_SP7nc0_line3, M7_GSP10_line0);
inv M7_GSP10_SP7nc1_Xo0(LocalCarryXCin0_25, M7_GSP10_SP7nc1_NotA);
inv M7_GSP10_SP7nc1_Xo1(M7_GSP10_line0, M7_GSP10_SP7nc1_NotB);
nand2 M7_GSP10_SP7nc1_Xo2(M7_GSP10_SP7nc1_NotA, M7_GSP10_line0, M7_GSP10_SP7nc1_line2);
nand2 M7_GSP10_SP7nc1_Xo3(M7_GSP10_SP7nc1_NotB, LocalCarryXCin0_25, M7_GSP10_SP7nc1_line3);
nand2 M7_GSP10_SP7nc1_Xo4(M7_GSP10_SP7nc1_line2, M7_GSP10_SP7nc1_line3, M7_GSP10_line1);
inv M7_GSP10_SP7nc2_Xo0(PropXbus_23, M7_GSP10_SP7nc2_NotA);
inv M7_GSP10_SP7nc2_Xo1(M7_GSP10_line1, M7_GSP10_SP7nc2_NotB);
nand2 M7_GSP10_SP7nc2_Xo2(M7_GSP10_SP7nc2_NotA, M7_GSP10_line1, M7_GSP10_SP7nc2_line2);
nand2 M7_GSP10_SP7nc2_Xo3(M7_GSP10_SP7nc2_NotB, PropXbus_23, M7_GSP10_SP7nc2_line3);
nand2 M7_GSP10_SP7nc2_Xo4(M7_GSP10_SP7nc2_line2, M7_GSP10_SP7nc2_line3, M7_GSP10_line2);
inv M7_GSP10_SP7nc3_Xo0(PropXbus_24, M7_GSP10_SP7nc3_NotA);
inv M7_GSP10_SP7nc3_Xo1(M7_GSP10_line2, M7_GSP10_SP7nc3_NotB);
nand2 M7_GSP10_SP7nc3_Xo2(M7_GSP10_SP7nc3_NotA, M7_GSP10_line2, M7_GSP10_SP7nc3_line2);
nand2 M7_GSP10_SP7nc3_Xo3(M7_GSP10_SP7nc3_NotB, PropXbus_24, M7_GSP10_SP7nc3_line3);
nand2 M7_GSP10_SP7nc3_Xo4(M7_GSP10_SP7nc3_line2, M7_GSP10_SP7nc3_line3, M7_GSP10_line3);
inv M7_GSP10_SP7nc4_Xo0(PropXbus_25, M7_GSP10_SP7nc4_NotA);
inv M7_GSP10_SP7nc4_Xo1(M7_GSP10_line3, M7_GSP10_SP7nc4_NotB);
nand2 M7_GSP10_SP7nc4_Xo2(M7_GSP10_SP7nc4_NotA, M7_GSP10_line3, M7_GSP10_SP7nc4_line2);
nand2 M7_GSP10_SP7nc4_Xo3(M7_GSP10_SP7nc4_NotB, PropXbus_25, M7_GSP10_SP7nc4_line3);
nand2 M7_GSP10_SP7nc4_Xo4(M7_GSP10_SP7nc4_line2, M7_GSP10_SP7nc4_line3, M7_GSP10_line4);
inv M7_GSP10_SP7nc5_Xo0(PropXbus_26, M7_GSP10_SP7nc5_NotA);
inv M7_GSP10_SP7nc5_Xo1(M7_GSP10_line4, M7_GSP10_SP7nc5_NotB);
nand2 M7_GSP10_SP7nc5_Xo2(M7_GSP10_SP7nc5_NotA, M7_GSP10_line4, M7_GSP10_SP7nc5_line2);
nand2 M7_GSP10_SP7nc5_Xo3(M7_GSP10_SP7nc5_NotB, PropXbus_26, M7_GSP10_SP7nc5_line3);
nand2 M7_GSP10_SP7nc5_Xo4(M7_GSP10_SP7nc5_line2, M7_GSP10_SP7nc5_line3, M7_ParCin0b26_23);
inv M7_GSP11_SP7c0(PropXbus_26, M7_GSP11_NewInbus_6);
inv M7_GSP11_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_23, M7_GSP11_SP7c2_SP7nc0_NotA);
inv M7_GSP11_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_24, M7_GSP11_SP7c2_SP7nc0_NotB);
nand2 M7_GSP11_SP7c2_SP7nc0_Xo2(M7_GSP11_SP7c2_SP7nc0_NotA, LocalCarryXCin1_24, M7_GSP11_SP7c2_SP7nc0_line2);
nand2 M7_GSP11_SP7c2_SP7nc0_Xo3(M7_GSP11_SP7c2_SP7nc0_NotB, LocalCarryXCin1_23, M7_GSP11_SP7c2_SP7nc0_line3);
nand2 M7_GSP11_SP7c2_SP7nc0_Xo4(M7_GSP11_SP7c2_SP7nc0_line2, M7_GSP11_SP7c2_SP7nc0_line3, M7_GSP11_SP7c2_line0);
inv M7_GSP11_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_25, M7_GSP11_SP7c2_SP7nc1_NotA);
inv M7_GSP11_SP7c2_SP7nc1_Xo1(M7_GSP11_SP7c2_line0, M7_GSP11_SP7c2_SP7nc1_NotB);
nand2 M7_GSP11_SP7c2_SP7nc1_Xo2(M7_GSP11_SP7c2_SP7nc1_NotA, M7_GSP11_SP7c2_line0, M7_GSP11_SP7c2_SP7nc1_line2);
nand2 M7_GSP11_SP7c2_SP7nc1_Xo3(M7_GSP11_SP7c2_SP7nc1_NotB, LocalCarryXCin1_25, M7_GSP11_SP7c2_SP7nc1_line3);
nand2 M7_GSP11_SP7c2_SP7nc1_Xo4(M7_GSP11_SP7c2_SP7nc1_line2, M7_GSP11_SP7c2_SP7nc1_line3, M7_GSP11_SP7c2_line1);
inv M7_GSP11_SP7c2_SP7nc2_Xo0(PropXbus_23, M7_GSP11_SP7c2_SP7nc2_NotA);
inv M7_GSP11_SP7c2_SP7nc2_Xo1(M7_GSP11_SP7c2_line1, M7_GSP11_SP7c2_SP7nc2_NotB);
nand2 M7_GSP11_SP7c2_SP7nc2_Xo2(M7_GSP11_SP7c2_SP7nc2_NotA, M7_GSP11_SP7c2_line1, M7_GSP11_SP7c2_SP7nc2_line2);
nand2 M7_GSP11_SP7c2_SP7nc2_Xo3(M7_GSP11_SP7c2_SP7nc2_NotB, PropXbus_23, M7_GSP11_SP7c2_SP7nc2_line3);
nand2 M7_GSP11_SP7c2_SP7nc2_Xo4(M7_GSP11_SP7c2_SP7nc2_line2, M7_GSP11_SP7c2_SP7nc2_line3, M7_GSP11_SP7c2_line2);
inv M7_GSP11_SP7c2_SP7nc3_Xo0(PropXbus_24, M7_GSP11_SP7c2_SP7nc3_NotA);
inv M7_GSP11_SP7c2_SP7nc3_Xo1(M7_GSP11_SP7c2_line2, M7_GSP11_SP7c2_SP7nc3_NotB);
nand2 M7_GSP11_SP7c2_SP7nc3_Xo2(M7_GSP11_SP7c2_SP7nc3_NotA, M7_GSP11_SP7c2_line2, M7_GSP11_SP7c2_SP7nc3_line2);
nand2 M7_GSP11_SP7c2_SP7nc3_Xo3(M7_GSP11_SP7c2_SP7nc3_NotB, PropXbus_24, M7_GSP11_SP7c2_SP7nc3_line3);
nand2 M7_GSP11_SP7c2_SP7nc3_Xo4(M7_GSP11_SP7c2_SP7nc3_line2, M7_GSP11_SP7c2_SP7nc3_line3, M7_GSP11_SP7c2_line3);
inv M7_GSP11_SP7c2_SP7nc4_Xo0(PropXbus_25, M7_GSP11_SP7c2_SP7nc4_NotA);
inv M7_GSP11_SP7c2_SP7nc4_Xo1(M7_GSP11_SP7c2_line3, M7_GSP11_SP7c2_SP7nc4_NotB);
nand2 M7_GSP11_SP7c2_SP7nc4_Xo2(M7_GSP11_SP7c2_SP7nc4_NotA, M7_GSP11_SP7c2_line3, M7_GSP11_SP7c2_SP7nc4_line2);
nand2 M7_GSP11_SP7c2_SP7nc4_Xo3(M7_GSP11_SP7c2_SP7nc4_NotB, PropXbus_25, M7_GSP11_SP7c2_SP7nc4_line3);
nand2 M7_GSP11_SP7c2_SP7nc4_Xo4(M7_GSP11_SP7c2_SP7nc4_line2, M7_GSP11_SP7c2_SP7nc4_line3, M7_GSP11_SP7c2_line4);
inv M7_GSP11_SP7c2_SP7nc5_Xo0(M7_GSP11_NewInbus_6, M7_GSP11_SP7c2_SP7nc5_NotA);
inv M7_GSP11_SP7c2_SP7nc5_Xo1(M7_GSP11_SP7c2_line4, M7_GSP11_SP7c2_SP7nc5_NotB);
nand2 M7_GSP11_SP7c2_SP7nc5_Xo2(M7_GSP11_SP7c2_SP7nc5_NotA, M7_GSP11_SP7c2_line4, M7_GSP11_SP7c2_SP7nc5_line2);
nand2 M7_GSP11_SP7c2_SP7nc5_Xo3(M7_GSP11_SP7c2_SP7nc5_NotB, M7_GSP11_NewInbus_6, M7_GSP11_SP7c2_SP7nc5_line3);
nand2 M7_GSP11_SP7c2_SP7nc5_Xo4(M7_GSP11_SP7c2_SP7nc5_line2, M7_GSP11_SP7c2_SP7nc5_line3, M7_ParCin1b26_23);
inv M7_GSP12_SP9nc0_SP7nc0_Xo0(M5_GenXbus_27, M7_GSP12_SP9nc0_SP7nc0_NotA);
inv M7_GSP12_SP9nc0_SP7nc0_Xo1(LocalCarryXCin0_28, M7_GSP12_SP9nc0_SP7nc0_NotB);
nand2 M7_GSP12_SP9nc0_SP7nc0_Xo2(M7_GSP12_SP9nc0_SP7nc0_NotA, LocalCarryXCin0_28, M7_GSP12_SP9nc0_SP7nc0_line2);
nand2 M7_GSP12_SP9nc0_SP7nc0_Xo3(M7_GSP12_SP9nc0_SP7nc0_NotB, M5_GenXbus_27, M7_GSP12_SP9nc0_SP7nc0_line3);
nand2 M7_GSP12_SP9nc0_SP7nc0_Xo4(M7_GSP12_SP9nc0_SP7nc0_line2, M7_GSP12_SP9nc0_SP7nc0_line3, M7_GSP12_SP9nc0_line0);
inv M7_GSP12_SP9nc0_SP7nc1_Xo0(LocalCarryXCin0_29, M7_GSP12_SP9nc0_SP7nc1_NotA);
inv M7_GSP12_SP9nc0_SP7nc1_Xo1(M7_GSP12_SP9nc0_line0, M7_GSP12_SP9nc0_SP7nc1_NotB);
nand2 M7_GSP12_SP9nc0_SP7nc1_Xo2(M7_GSP12_SP9nc0_SP7nc1_NotA, M7_GSP12_SP9nc0_line0, M7_GSP12_SP9nc0_SP7nc1_line2);
nand2 M7_GSP12_SP9nc0_SP7nc1_Xo3(M7_GSP12_SP9nc0_SP7nc1_NotB, LocalCarryXCin0_29, M7_GSP12_SP9nc0_SP7nc1_line3);
nand2 M7_GSP12_SP9nc0_SP7nc1_Xo4(M7_GSP12_SP9nc0_SP7nc1_line2, M7_GSP12_SP9nc0_SP7nc1_line3, M7_GSP12_SP9nc0_line1);
inv M7_GSP12_SP9nc0_SP7nc2_Xo0(LocalCarryXCin0_30, M7_GSP12_SP9nc0_SP7nc2_NotA);
inv M7_GSP12_SP9nc0_SP7nc2_Xo1(M7_GSP12_SP9nc0_line1, M7_GSP12_SP9nc0_SP7nc2_NotB);
nand2 M7_GSP12_SP9nc0_SP7nc2_Xo2(M7_GSP12_SP9nc0_SP7nc2_NotA, M7_GSP12_SP9nc0_line1, M7_GSP12_SP9nc0_SP7nc2_line2);
nand2 M7_GSP12_SP9nc0_SP7nc2_Xo3(M7_GSP12_SP9nc0_SP7nc2_NotB, LocalCarryXCin0_30, M7_GSP12_SP9nc0_SP7nc2_line3);
nand2 M7_GSP12_SP9nc0_SP7nc2_Xo4(M7_GSP12_SP9nc0_SP7nc2_line2, M7_GSP12_SP9nc0_SP7nc2_line3, M7_GSP12_SP9nc0_line2);
inv M7_GSP12_SP9nc0_SP7nc3_Xo0(PropXbus_27, M7_GSP12_SP9nc0_SP7nc3_NotA);
inv M7_GSP12_SP9nc0_SP7nc3_Xo1(M7_GSP12_SP9nc0_line2, M7_GSP12_SP9nc0_SP7nc3_NotB);
nand2 M7_GSP12_SP9nc0_SP7nc3_Xo2(M7_GSP12_SP9nc0_SP7nc3_NotA, M7_GSP12_SP9nc0_line2, M7_GSP12_SP9nc0_SP7nc3_line2);
nand2 M7_GSP12_SP9nc0_SP7nc3_Xo3(M7_GSP12_SP9nc0_SP7nc3_NotB, PropXbus_27, M7_GSP12_SP9nc0_SP7nc3_line3);
nand2 M7_GSP12_SP9nc0_SP7nc3_Xo4(M7_GSP12_SP9nc0_SP7nc3_line2, M7_GSP12_SP9nc0_SP7nc3_line3, M7_GSP12_SP9nc0_line3);
inv M7_GSP12_SP9nc0_SP7nc4_Xo0(PropXbus_28, M7_GSP12_SP9nc0_SP7nc4_NotA);
inv M7_GSP12_SP9nc0_SP7nc4_Xo1(M7_GSP12_SP9nc0_line3, M7_GSP12_SP9nc0_SP7nc4_NotB);
nand2 M7_GSP12_SP9nc0_SP7nc4_Xo2(M7_GSP12_SP9nc0_SP7nc4_NotA, M7_GSP12_SP9nc0_line3, M7_GSP12_SP9nc0_SP7nc4_line2);
nand2 M7_GSP12_SP9nc0_SP7nc4_Xo3(M7_GSP12_SP9nc0_SP7nc4_NotB, PropXbus_28, M7_GSP12_SP9nc0_SP7nc4_line3);
nand2 M7_GSP12_SP9nc0_SP7nc4_Xo4(M7_GSP12_SP9nc0_SP7nc4_line2, M7_GSP12_SP9nc0_SP7nc4_line3, M7_GSP12_SP9nc0_line4);
inv M7_GSP12_SP9nc0_SP7nc5_Xo0(PropXbus_29, M7_GSP12_SP9nc0_SP7nc5_NotA);
inv M7_GSP12_SP9nc0_SP7nc5_Xo1(M7_GSP12_SP9nc0_line4, M7_GSP12_SP9nc0_SP7nc5_NotB);
nand2 M7_GSP12_SP9nc0_SP7nc5_Xo2(M7_GSP12_SP9nc0_SP7nc5_NotA, M7_GSP12_SP9nc0_line4, M7_GSP12_SP9nc0_SP7nc5_line2);
nand2 M7_GSP12_SP9nc0_SP7nc5_Xo3(M7_GSP12_SP9nc0_SP7nc5_NotB, PropXbus_29, M7_GSP12_SP9nc0_SP7nc5_line3);
nand2 M7_GSP12_SP9nc0_SP7nc5_Xo4(M7_GSP12_SP9nc0_SP7nc5_line2, M7_GSP12_SP9nc0_SP7nc5_line3, M7_GSP12_line0);
inv M7_GSP12_SP9nc1_Xo0(PropXbus_30, M7_GSP12_SP9nc1_NotA);
inv M7_GSP12_SP9nc1_Xo1(M7_GSP12_line0, M7_GSP12_SP9nc1_NotB);
nand2 M7_GSP12_SP9nc1_Xo2(M7_GSP12_SP9nc1_NotA, M7_GSP12_line0, M7_GSP12_SP9nc1_line2);
nand2 M7_GSP12_SP9nc1_Xo3(M7_GSP12_SP9nc1_NotB, PropXbus_30, M7_GSP12_SP9nc1_line3);
nand2 M7_GSP12_SP9nc1_Xo4(M7_GSP12_SP9nc1_line2, M7_GSP12_SP9nc1_line3, M7_GSP12_line1);
inv M7_GSP12_SP9nc2_Xo0(PropXbus_31, M7_GSP12_SP9nc2_NotA);
inv M7_GSP12_SP9nc2_Xo1(M7_GSP12_line1, M7_GSP12_SP9nc2_NotB);
nand2 M7_GSP12_SP9nc2_Xo2(M7_GSP12_SP9nc2_NotA, M7_GSP12_line1, M7_GSP12_SP9nc2_line2);
nand2 M7_GSP12_SP9nc2_Xo3(M7_GSP12_SP9nc2_NotB, PropXbus_31, M7_GSP12_SP9nc2_line3);
nand2 M7_GSP12_SP9nc2_Xo4(M7_GSP12_SP9nc2_line2, M7_GSP12_SP9nc2_line3, M7_ParCin0b31_27);
inv M7_GSP13_SP9nc0_SP7c0(PropXbus_29, M7_GSP13_SP9nc0_NewInbus_6);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc0_Xo0(LocalCarryXCin1_27, M7_GSP13_SP9nc0_SP7c2_SP7nc0_NotA);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc0_Xo1(LocalCarryXCin1_28, M7_GSP13_SP9nc0_SP7c2_SP7nc0_NotB);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc0_Xo2(M7_GSP13_SP9nc0_SP7c2_SP7nc0_NotA, LocalCarryXCin1_28, M7_GSP13_SP9nc0_SP7c2_SP7nc0_line2);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc0_Xo3(M7_GSP13_SP9nc0_SP7c2_SP7nc0_NotB, LocalCarryXCin1_27, M7_GSP13_SP9nc0_SP7c2_SP7nc0_line3);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc0_Xo4(M7_GSP13_SP9nc0_SP7c2_SP7nc0_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc0_line3, M7_GSP13_SP9nc0_SP7c2_line0);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc1_Xo0(LocalCarryXCin1_29, M7_GSP13_SP9nc0_SP7c2_SP7nc1_NotA);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc1_Xo1(M7_GSP13_SP9nc0_SP7c2_line0, M7_GSP13_SP9nc0_SP7c2_SP7nc1_NotB);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc1_Xo2(M7_GSP13_SP9nc0_SP7c2_SP7nc1_NotA, M7_GSP13_SP9nc0_SP7c2_line0, M7_GSP13_SP9nc0_SP7c2_SP7nc1_line2);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc1_Xo3(M7_GSP13_SP9nc0_SP7c2_SP7nc1_NotB, LocalCarryXCin1_29, M7_GSP13_SP9nc0_SP7c2_SP7nc1_line3);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc1_Xo4(M7_GSP13_SP9nc0_SP7c2_SP7nc1_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc1_line3, M7_GSP13_SP9nc0_SP7c2_line1);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc2_Xo0(LocalCarryXCin1_30, M7_GSP13_SP9nc0_SP7c2_SP7nc2_NotA);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc2_Xo1(M7_GSP13_SP9nc0_SP7c2_line1, M7_GSP13_SP9nc0_SP7c2_SP7nc2_NotB);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc2_Xo2(M7_GSP13_SP9nc0_SP7c2_SP7nc2_NotA, M7_GSP13_SP9nc0_SP7c2_line1, M7_GSP13_SP9nc0_SP7c2_SP7nc2_line2);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc2_Xo3(M7_GSP13_SP9nc0_SP7c2_SP7nc2_NotB, LocalCarryXCin1_30, M7_GSP13_SP9nc0_SP7c2_SP7nc2_line3);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc2_Xo4(M7_GSP13_SP9nc0_SP7c2_SP7nc2_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc2_line3, M7_GSP13_SP9nc0_SP7c2_line2);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc3_Xo0(PropXbus_27, M7_GSP13_SP9nc0_SP7c2_SP7nc3_NotA);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc3_Xo1(M7_GSP13_SP9nc0_SP7c2_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc3_NotB);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc3_Xo2(M7_GSP13_SP9nc0_SP7c2_SP7nc3_NotA, M7_GSP13_SP9nc0_SP7c2_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc3_line2);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc3_Xo3(M7_GSP13_SP9nc0_SP7c2_SP7nc3_NotB, PropXbus_27, M7_GSP13_SP9nc0_SP7c2_SP7nc3_line3);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc3_Xo4(M7_GSP13_SP9nc0_SP7c2_SP7nc3_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc3_line3, M7_GSP13_SP9nc0_SP7c2_line3);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc4_Xo0(PropXbus_28, M7_GSP13_SP9nc0_SP7c2_SP7nc4_NotA);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc4_Xo1(M7_GSP13_SP9nc0_SP7c2_line3, M7_GSP13_SP9nc0_SP7c2_SP7nc4_NotB);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc4_Xo2(M7_GSP13_SP9nc0_SP7c2_SP7nc4_NotA, M7_GSP13_SP9nc0_SP7c2_line3, M7_GSP13_SP9nc0_SP7c2_SP7nc4_line2);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc4_Xo3(M7_GSP13_SP9nc0_SP7c2_SP7nc4_NotB, PropXbus_28, M7_GSP13_SP9nc0_SP7c2_SP7nc4_line3);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc4_Xo4(M7_GSP13_SP9nc0_SP7c2_SP7nc4_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc4_line3, M7_GSP13_SP9nc0_SP7c2_line4);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc5_Xo0(M7_GSP13_SP9nc0_NewInbus_6, M7_GSP13_SP9nc0_SP7c2_SP7nc5_NotA);
inv M7_GSP13_SP9nc0_SP7c2_SP7nc5_Xo1(M7_GSP13_SP9nc0_SP7c2_line4, M7_GSP13_SP9nc0_SP7c2_SP7nc5_NotB);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc5_Xo2(M7_GSP13_SP9nc0_SP7c2_SP7nc5_NotA, M7_GSP13_SP9nc0_SP7c2_line4, M7_GSP13_SP9nc0_SP7c2_SP7nc5_line2);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc5_Xo3(M7_GSP13_SP9nc0_SP7c2_SP7nc5_NotB, M7_GSP13_SP9nc0_NewInbus_6, M7_GSP13_SP9nc0_SP7c2_SP7nc5_line3);
nand2 M7_GSP13_SP9nc0_SP7c2_SP7nc5_Xo4(M7_GSP13_SP9nc0_SP7c2_SP7nc5_line2, M7_GSP13_SP9nc0_SP7c2_SP7nc5_line3, M7_GSP13_line0);
inv M7_GSP13_SP9nc1_Xo0(PropXbus_30, M7_GSP13_SP9nc1_NotA);
inv M7_GSP13_SP9nc1_Xo1(M7_GSP13_line0, M7_GSP13_SP9nc1_NotB);
nand2 M7_GSP13_SP9nc1_Xo2(M7_GSP13_SP9nc1_NotA, M7_GSP13_line0, M7_GSP13_SP9nc1_line2);
nand2 M7_GSP13_SP9nc1_Xo3(M7_GSP13_SP9nc1_NotB, PropXbus_30, M7_GSP13_SP9nc1_line3);
nand2 M7_GSP13_SP9nc1_Xo4(M7_GSP13_SP9nc1_line2, M7_GSP13_SP9nc1_line3, M7_GSP13_line1);
inv M7_GSP13_SP9nc2_Xo0(PropXbus_31, M7_GSP13_SP9nc2_NotA);
inv M7_GSP13_SP9nc2_Xo1(M7_GSP13_line1, M7_GSP13_SP9nc2_NotB);
nand2 M7_GSP13_SP9nc2_Xo2(M7_GSP13_SP9nc2_NotA, M7_GSP13_line1, M7_GSP13_SP9nc2_line2);
nand2 M7_GSP13_SP9nc2_Xo3(M7_GSP13_SP9nc2_NotB, PropXbus_31, M7_GSP13_SP9nc2_line3);
nand2 M7_GSP13_SP9nc2_Xo4(M7_GSP13_SP9nc2_line2, M7_GSP13_SP9nc2_line3, M7_ParCin1b31_27);
inv M7_GSP14_SP3nc0_Xo0(M5_GenXbus_32, M7_GSP14_SP3nc0_NotA);
inv M7_GSP14_SP3nc0_Xo1(PropXbus_32, M7_GSP14_SP3nc0_NotB);
nand2 M7_GSP14_SP3nc0_Xo2(M7_GSP14_SP3nc0_NotA, PropXbus_32, M7_GSP14_SP3nc0_line2);
nand2 M7_GSP14_SP3nc0_Xo3(M7_GSP14_SP3nc0_NotB, M5_GenXbus_32, M7_GSP14_SP3nc0_line3);
nand2 M7_GSP14_SP3nc0_Xo4(M7_GSP14_SP3nc0_line2, M7_GSP14_SP3nc0_line3, M7_GSP14_line0);
inv M7_GSP14_SP3nc1_Xo0(PropXbus_33, M7_GSP14_SP3nc1_NotA);
inv M7_GSP14_SP3nc1_Xo1(M7_GSP14_line0, M7_GSP14_SP3nc1_NotB);
nand2 M7_GSP14_SP3nc1_Xo2(M7_GSP14_SP3nc1_NotA, M7_GSP14_line0, M7_GSP14_SP3nc1_line2);
nand2 M7_GSP14_SP3nc1_Xo3(M7_GSP14_SP3nc1_NotB, PropXbus_33, M7_GSP14_SP3nc1_line3);
nand2 M7_GSP14_SP3nc1_Xo4(M7_GSP14_SP3nc1_line2, M7_GSP14_SP3nc1_line3, M7_ParCin0b33_32);
inv M7_GSP15_SP3c0(PropXbus_33, M7_GSP15_NotIn2);
inv M7_GSP15_SP3c1_Xo0(LocalCarryXCin1_32, M7_GSP15_SP3c1_NotA);
inv M7_GSP15_SP3c1_Xo1(PropXbus_32, M7_GSP15_SP3c1_NotB);
nand2 M7_GSP15_SP3c1_Xo2(M7_GSP15_SP3c1_NotA, PropXbus_32, M7_GSP15_SP3c1_line2);
nand2 M7_GSP15_SP3c1_Xo3(M7_GSP15_SP3c1_NotB, LocalCarryXCin1_32, M7_GSP15_SP3c1_line3);
nand2 M7_GSP15_SP3c1_Xo4(M7_GSP15_SP3c1_line2, M7_GSP15_SP3c1_line3, M7_GSP15_line1);
inv M7_GSP15_SP3c2_Xo0(M7_GSP15_NotIn2, M7_GSP15_SP3c2_NotA);
inv M7_GSP15_SP3c2_Xo1(M7_GSP15_line1, M7_GSP15_SP3c2_NotB);
nand2 M7_GSP15_SP3c2_Xo2(M7_GSP15_SP3c2_NotA, M7_GSP15_line1, M7_GSP15_SP3c2_line2);
nand2 M7_GSP15_SP3c2_Xo3(M7_GSP15_SP3c2_NotB, M7_GSP15_NotIn2, M7_GSP15_SP3c2_line3);
nand2 M7_GSP15_SP3c2_Xo4(M7_GSP15_SP3c2_line2, M7_GSP15_SP3c2_line3, M7_ParCin1b33_32armut);
inv M7_GSP16_SPar0_Mux0(in4526, M7_GSP16_SPar0_Not_ContIn);
and2 M7_GSP16_SPar0_Mux1(M7_ParCin0b4_0, M7_GSP16_SPar0_Not_ContIn, M7_GSP16_SPar0_line1);
and2 M7_GSP16_SPar0_Mux2(M7_ParCin1b4_0, in4526, M7_GSP16_SPar0_line2);
or2 M7_GSP16_SPar0_Mux3(M7_GSP16_SPar0_line1, M7_GSP16_SPar0_line2, M7_GSP16_line0);
inv M7_GSP16_SPar1_Mux0(LocalCarryXCin0_4, M7_GSP16_SPar1_Not_ContIn);
and2 M7_GSP16_SPar1_Mux1(M7_ParCin0b8_5, M7_GSP16_SPar1_Not_ContIn, M7_GSP16_SPar1_line1);
and2 M7_GSP16_SPar1_Mux2(M7_ParCin1b8_5, LocalCarryXCin0_4, M7_GSP16_SPar1_line2);
or2 M7_GSP16_SPar1_Mux3(M7_GSP16_SPar1_line1, M7_GSP16_SPar1_line2, M7_GSP16_line1);
inv M7_GSP16_SPar2_Mux0(LocalCarryXCin1_4, M7_GSP16_SPar2_Not_ContIn);
and2 M7_GSP16_SPar2_Mux1(M7_ParCin0b8_5, M7_GSP16_SPar2_Not_ContIn, M7_GSP16_SPar2_line1);
and2 M7_GSP16_SPar2_Mux2(M7_ParCin1b8_5, LocalCarryXCin1_4, M7_GSP16_SPar2_line2);
or2 M7_GSP16_SPar2_Mux3(M7_GSP16_SPar2_line1, M7_GSP16_SPar2_line2, M7_GSP16_line2);
inv M7_GSP16_SPar3_Mux0(in4526, M7_GSP16_SPar3_Not_ContIn);
and2 M7_GSP16_SPar3_Mux1(M7_GSP16_line1, M7_GSP16_SPar3_Not_ContIn, M7_GSP16_SPar3_line1);
and2 M7_GSP16_SPar3_Mux2(M7_GSP16_line2, in4526, M7_GSP16_SPar3_line2);
or2 M7_GSP16_SPar3_Mux3(M7_GSP16_SPar3_line1, M7_GSP16_SPar3_line2, M7_GSP16_line3);
inv M7_GSP16_SPar4_Xo0(M7_GSP16_line0, M7_GSP16_SPar4_NotA);
inv M7_GSP16_SPar4_Xo1(M7_GSP16_line3, M7_GSP16_SPar4_NotB);
nand2 M7_GSP16_SPar4_Xo2(M7_GSP16_SPar4_NotA, M7_GSP16_line3, M7_GSP16_SPar4_line2);
nand2 M7_GSP16_SPar4_Xo3(M7_GSP16_SPar4_NotB, M7_GSP16_line0, M7_GSP16_SPar4_line3);
nand2 M7_GSP16_SPar4_Xo4(M7_GSP16_SPar4_line2, M7_GSP16_SPar4_line3, M7_GSP16_line4);
inv M7_GSP16_SPar5(M7_GSP16_line4, out399);
inv M7_GSP17_SPar0_Mux0(CarryXbus_8, M7_GSP17_SPar0_Not_ContIn);
and2 M7_GSP17_SPar0_Mux1(M7_ParCin0b13_9, M7_GSP17_SPar0_Not_ContIn, M7_GSP17_SPar0_line1);
and2 M7_GSP17_SPar0_Mux2(M7_ParCin1b13_9, CarryXbus_8, M7_GSP17_SPar0_line2);
or2 M7_GSP17_SPar0_Mux3(M7_GSP17_SPar0_line1, M7_GSP17_SPar0_line2, M7_GSP17_line0);
inv M7_GSP17_SPar1_Mux0(LocalCarryXCin0_13, M7_GSP17_SPar1_Not_ContIn);
and2 M7_GSP17_SPar1_Mux1(M7_ParCin0b17_14, M7_GSP17_SPar1_Not_ContIn, M7_GSP17_SPar1_line1);
and2 M7_GSP17_SPar1_Mux2(M7_ParCin1b17_14, LocalCarryXCin0_13, M7_GSP17_SPar1_line2);
or2 M7_GSP17_SPar1_Mux3(M7_GSP17_SPar1_line1, M7_GSP17_SPar1_line2, M7_GSP17_line1);
inv M7_GSP17_SPar2_Mux0(LocalCarryXCin1_13, M7_GSP17_SPar2_Not_ContIn);
and2 M7_GSP17_SPar2_Mux1(M7_ParCin0b17_14, M7_GSP17_SPar2_Not_ContIn, M7_GSP17_SPar2_line1);
and2 M7_GSP17_SPar2_Mux2(M7_ParCin1b17_14, LocalCarryXCin1_13, M7_GSP17_SPar2_line2);
or2 M7_GSP17_SPar2_Mux3(M7_GSP17_SPar2_line1, M7_GSP17_SPar2_line2, M7_GSP17_line2);
inv M7_GSP17_SPar3_Mux0(CarryXbus_8, M7_GSP17_SPar3_Not_ContIn);
and2 M7_GSP17_SPar3_Mux1(M7_GSP17_line1, M7_GSP17_SPar3_Not_ContIn, M7_GSP17_SPar3_line1);
and2 M7_GSP17_SPar3_Mux2(M7_GSP17_line2, CarryXbus_8, M7_GSP17_SPar3_line2);
or2 M7_GSP17_SPar3_Mux3(M7_GSP17_SPar3_line1, M7_GSP17_SPar3_line2, M7_GSP17_line3);
inv M7_GSP17_SPar4_Xo0(M7_GSP17_line0, M7_GSP17_SPar4_NotA);
inv M7_GSP17_SPar4_Xo1(M7_GSP17_line3, M7_GSP17_SPar4_NotB);
nand2 M7_GSP17_SPar4_Xo2(M7_GSP17_SPar4_NotA, M7_GSP17_line3, M7_GSP17_SPar4_line2);
nand2 M7_GSP17_SPar4_Xo3(M7_GSP17_SPar4_NotB, M7_GSP17_line0, M7_GSP17_SPar4_line3);
nand2 M7_GSP17_SPar4_Xo4(M7_GSP17_SPar4_line2, M7_GSP17_SPar4_line3, M7_GSP17_line4);
inv M7_GSP17_SPar5(M7_GSP17_line4, out370);
inv M7_GSP18_SPar0_Mux0(CarryXbus_17, M7_GSP18_SPar0_Not_ContIn);
and2 M7_GSP18_SPar0_Mux1(M7_ParCin0b22_18, M7_GSP18_SPar0_Not_ContIn, M7_GSP18_SPar0_line1);
and2 M7_GSP18_SPar0_Mux2(M7_ParCin1b22_18, CarryXbus_17, M7_GSP18_SPar0_line2);
or2 M7_GSP18_SPar0_Mux3(M7_GSP18_SPar0_line1, M7_GSP18_SPar0_line2, M7_GSP18_line0);
inv M7_GSP18_SPar1_Mux0(LocalCarryXCin0_22, M7_GSP18_SPar1_Not_ContIn);
and2 M7_GSP18_SPar1_Mux1(M7_ParCin0b26_23, M7_GSP18_SPar1_Not_ContIn, M7_GSP18_SPar1_line1);
and2 M7_GSP18_SPar1_Mux2(M7_ParCin1b26_23, LocalCarryXCin0_22, M7_GSP18_SPar1_line2);
or2 M7_GSP18_SPar1_Mux3(M7_GSP18_SPar1_line1, M7_GSP18_SPar1_line2, M7_GSP18_line1);
inv M7_GSP18_SPar2_Mux0(LocalCarryXCin1_22, M7_GSP18_SPar2_Not_ContIn);
and2 M7_GSP18_SPar2_Mux1(M7_ParCin0b26_23, M7_GSP18_SPar2_Not_ContIn, M7_GSP18_SPar2_line1);
and2 M7_GSP18_SPar2_Mux2(M7_ParCin1b26_23, LocalCarryXCin1_22, M7_GSP18_SPar2_line2);
or2 M7_GSP18_SPar2_Mux3(M7_GSP18_SPar2_line1, M7_GSP18_SPar2_line2, M7_GSP18_line2);
inv M7_GSP18_SPar3_Mux0(CarryXbus_17, M7_GSP18_SPar3_Not_ContIn);
and2 M7_GSP18_SPar3_Mux1(M7_GSP18_line1, M7_GSP18_SPar3_Not_ContIn, M7_GSP18_SPar3_line1);
and2 M7_GSP18_SPar3_Mux2(M7_GSP18_line2, CarryXbus_17, M7_GSP18_SPar3_line2);
or2 M7_GSP18_SPar3_Mux3(M7_GSP18_SPar3_line1, M7_GSP18_SPar3_line2, M7_GSP18_line3);
inv M7_GSP18_SPar4_Xo0(M7_GSP18_line0, M7_GSP18_SPar4_NotA);
inv M7_GSP18_SPar4_Xo1(M7_GSP18_line3, M7_GSP18_SPar4_NotB);
nand2 M7_GSP18_SPar4_Xo2(M7_GSP18_SPar4_NotA, M7_GSP18_line3, M7_GSP18_SPar4_line2);
nand2 M7_GSP18_SPar4_Xo3(M7_GSP18_SPar4_NotB, M7_GSP18_line0, M7_GSP18_SPar4_line3);
nand2 M7_GSP18_SPar4_Xo4(M7_GSP18_SPar4_line2, M7_GSP18_SPar4_line3, M7_GSP18_line4);
inv M7_GSP18_SPar5(M7_GSP18_line4, out321);
inv M7_GSP19_SPar0_Mux0(CarryXbus_26, M7_GSP19_SPar0_Not_ContIn);
and2 M7_GSP19_SPar0_Mux1(M7_ParCin0b31_27, M7_GSP19_SPar0_Not_ContIn, M7_GSP19_SPar0_line1);
and2 M7_GSP19_SPar0_Mux2(M7_ParCin1b31_27, CarryXbus_26, M7_GSP19_SPar0_line2);
or2 M7_GSP19_SPar0_Mux3(M7_GSP19_SPar0_line1, M7_GSP19_SPar0_line2, M7_GSP19_line0);
inv M7_GSP19_SPar1_Mux0(LocalCarryXCin0_31, M7_GSP19_SPar1_Not_ContIn);
and2 M7_GSP19_SPar1_Mux1(M7_ParCin0b33_32, M7_GSP19_SPar1_Not_ContIn, M7_GSP19_SPar1_line1);
and2 M7_GSP19_SPar1_Mux2(M7_ParCin1b33_32armut, LocalCarryXCin0_31, M7_GSP19_SPar1_line2);
or2 M7_GSP19_SPar1_Mux3(M7_GSP19_SPar1_line1, M7_GSP19_SPar1_line2, M7_GSP19_line1);
inv M7_GSP19_SPar2_Mux0(LocalCarryXCin1_31, M7_GSP19_SPar2_Not_ContIn);
and2 M7_GSP19_SPar2_Mux1(M7_ParCin0b33_32, M7_GSP19_SPar2_Not_ContIn, M7_GSP19_SPar2_line1);
and2 M7_GSP19_SPar2_Mux2(M7_ParCin1b33_32armut, LocalCarryXCin1_31, M7_GSP19_SPar2_line2);
or2 M7_GSP19_SPar2_Mux3(M7_GSP19_SPar2_line1, M7_GSP19_SPar2_line2, M7_GSP19_line2);
inv M7_GSP19_SPar3_Mux0(CarryXbus_26, M7_GSP19_SPar3_Not_ContIn);
and2 M7_GSP19_SPar3_Mux1(M7_GSP19_line1, M7_GSP19_SPar3_Not_ContIn, M7_GSP19_SPar3_line1);
and2 M7_GSP19_SPar3_Mux2(M7_GSP19_line2, CarryXbus_26, M7_GSP19_SPar3_line2);
or2 M7_GSP19_SPar3_Mux3(M7_GSP19_SPar3_line1, M7_GSP19_SPar3_line2, M7_GSP19_line3);
inv M7_GSP19_SPar4_Xo0(M7_GSP19_line0, M7_GSP19_SPar4_NotA);
inv M7_GSP19_SPar4_Xo1(M7_GSP19_line3, M7_GSP19_SPar4_NotB);
nand2 M7_GSP19_SPar4_Xo2(M7_GSP19_SPar4_NotA, M7_GSP19_line3, M7_GSP19_SPar4_line2);
nand2 M7_GSP19_SPar4_Xo3(M7_GSP19_SPar4_NotB, M7_GSP19_line0, M7_GSP19_SPar4_line3);
nand2 M7_GSP19_SPar4_Xo4(M7_GSP19_SPar4_line2, M7_GSP19_SPar4_line3, M7_GSP19_line4);
inv M7_GSP19_SPar5(M7_GSP19_line4, out338);
and2 M8_UM8_0_GP34_0_GenProp8_0(YAbus_0, YBbus_0, M8_GenYbus_0);
and2 M8_UM8_0_GP34_0_GenProp8_1(YAbus_1, YBbus_1, M8_GenYbus_1);
and2 M8_UM8_0_GP34_0_GenProp8_2(YAbus_2, YBbus_2, M8_GenYbus_2);
and2 M8_UM8_0_GP34_0_GenProp8_3(YAbus_3, YBbus_3, M8_GenYbus_3);
and2 M8_UM8_0_GP34_0_GenProp8_4(YAbus_4, YBbus_4, M8_GenYbus_4);
and2 M8_UM8_0_GP34_0_GenProp8_5(YAbus_5, YBbus_5, M8_GenYbus_5);
and2 M8_UM8_0_GP34_0_GenProp8_6(YAbus_6, YBbus_6, M8_GenYbus_6);
and2 M8_UM8_0_GP34_0_GenProp8_7(YAbus_7, YBbus_7, M8_GenYbus_7);
inv M8_UM8_0_GP34_0_GenProp8_8_Xo0(YAbus_0, M8_UM8_0_GP34_0_GenProp8_8_NotA);
inv M8_UM8_0_GP34_0_GenProp8_8_Xo1(YBbus_0, M8_UM8_0_GP34_0_GenProp8_8_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_8_Xo2(M8_UM8_0_GP34_0_GenProp8_8_NotA, YBbus_0, M8_UM8_0_GP34_0_GenProp8_8_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_8_Xo3(M8_UM8_0_GP34_0_GenProp8_8_NotB, YAbus_0, M8_UM8_0_GP34_0_GenProp8_8_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_8_Xo4(M8_UM8_0_GP34_0_GenProp8_8_line2, M8_UM8_0_GP34_0_GenProp8_8_line3, M8_PropYbus_0);
inv M8_UM8_0_GP34_0_GenProp8_9_Xo0(YAbus_1, M8_UM8_0_GP34_0_GenProp8_9_NotA);
inv M8_UM8_0_GP34_0_GenProp8_9_Xo1(YBbus_1, M8_UM8_0_GP34_0_GenProp8_9_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_9_Xo2(M8_UM8_0_GP34_0_GenProp8_9_NotA, YBbus_1, M8_UM8_0_GP34_0_GenProp8_9_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_9_Xo3(M8_UM8_0_GP34_0_GenProp8_9_NotB, YAbus_1, M8_UM8_0_GP34_0_GenProp8_9_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_9_Xo4(M8_UM8_0_GP34_0_GenProp8_9_line2, M8_UM8_0_GP34_0_GenProp8_9_line3, M8_PropYbus_1);
inv M8_UM8_0_GP34_0_GenProp8_10_Xo0(YAbus_2, M8_UM8_0_GP34_0_GenProp8_10_NotA);
inv M8_UM8_0_GP34_0_GenProp8_10_Xo1(YBbus_2, M8_UM8_0_GP34_0_GenProp8_10_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_10_Xo2(M8_UM8_0_GP34_0_GenProp8_10_NotA, YBbus_2, M8_UM8_0_GP34_0_GenProp8_10_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_10_Xo3(M8_UM8_0_GP34_0_GenProp8_10_NotB, YAbus_2, M8_UM8_0_GP34_0_GenProp8_10_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_10_Xo4(M8_UM8_0_GP34_0_GenProp8_10_line2, M8_UM8_0_GP34_0_GenProp8_10_line3, M8_PropYbus_2);
inv M8_UM8_0_GP34_0_GenProp8_11_Xo0(YAbus_3, M8_UM8_0_GP34_0_GenProp8_11_NotA);
inv M8_UM8_0_GP34_0_GenProp8_11_Xo1(YBbus_3, M8_UM8_0_GP34_0_GenProp8_11_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_11_Xo2(M8_UM8_0_GP34_0_GenProp8_11_NotA, YBbus_3, M8_UM8_0_GP34_0_GenProp8_11_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_11_Xo3(M8_UM8_0_GP34_0_GenProp8_11_NotB, YAbus_3, M8_UM8_0_GP34_0_GenProp8_11_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_11_Xo4(M8_UM8_0_GP34_0_GenProp8_11_line2, M8_UM8_0_GP34_0_GenProp8_11_line3, M8_PropYbus_3);
inv M8_UM8_0_GP34_0_GenProp8_12_Xo0(YAbus_4, M8_UM8_0_GP34_0_GenProp8_12_NotA);
inv M8_UM8_0_GP34_0_GenProp8_12_Xo1(YBbus_4, M8_UM8_0_GP34_0_GenProp8_12_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_12_Xo2(M8_UM8_0_GP34_0_GenProp8_12_NotA, YBbus_4, M8_UM8_0_GP34_0_GenProp8_12_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_12_Xo3(M8_UM8_0_GP34_0_GenProp8_12_NotB, YAbus_4, M8_UM8_0_GP34_0_GenProp8_12_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_12_Xo4(M8_UM8_0_GP34_0_GenProp8_12_line2, M8_UM8_0_GP34_0_GenProp8_12_line3, M8_PropYbus_4);
inv M8_UM8_0_GP34_0_GenProp8_13_Xo0(YAbus_5, M8_UM8_0_GP34_0_GenProp8_13_NotA);
inv M8_UM8_0_GP34_0_GenProp8_13_Xo1(YBbus_5, M8_UM8_0_GP34_0_GenProp8_13_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_13_Xo2(M8_UM8_0_GP34_0_GenProp8_13_NotA, YBbus_5, M8_UM8_0_GP34_0_GenProp8_13_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_13_Xo3(M8_UM8_0_GP34_0_GenProp8_13_NotB, YAbus_5, M8_UM8_0_GP34_0_GenProp8_13_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_13_Xo4(M8_UM8_0_GP34_0_GenProp8_13_line2, M8_UM8_0_GP34_0_GenProp8_13_line3, M8_PropYbus_5);
inv M8_UM8_0_GP34_0_GenProp8_14_Xo0(YAbus_6, M8_UM8_0_GP34_0_GenProp8_14_NotA);
inv M8_UM8_0_GP34_0_GenProp8_14_Xo1(YBbus_6, M8_UM8_0_GP34_0_GenProp8_14_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_14_Xo2(M8_UM8_0_GP34_0_GenProp8_14_NotA, YBbus_6, M8_UM8_0_GP34_0_GenProp8_14_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_14_Xo3(M8_UM8_0_GP34_0_GenProp8_14_NotB, YAbus_6, M8_UM8_0_GP34_0_GenProp8_14_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_14_Xo4(M8_UM8_0_GP34_0_GenProp8_14_line2, M8_UM8_0_GP34_0_GenProp8_14_line3, M8_PropYbus_6);
inv M8_UM8_0_GP34_0_GenProp8_15_Xo0(YAbus_7, M8_UM8_0_GP34_0_GenProp8_15_NotA);
inv M8_UM8_0_GP34_0_GenProp8_15_Xo1(YBbus_7, M8_UM8_0_GP34_0_GenProp8_15_NotB);
nand2 M8_UM8_0_GP34_0_GenProp8_15_Xo2(M8_UM8_0_GP34_0_GenProp8_15_NotA, YBbus_7, M8_UM8_0_GP34_0_GenProp8_15_line2);
nand2 M8_UM8_0_GP34_0_GenProp8_15_Xo3(M8_UM8_0_GP34_0_GenProp8_15_NotB, YAbus_7, M8_UM8_0_GP34_0_GenProp8_15_line3);
nand2 M8_UM8_0_GP34_0_GenProp8_15_Xo4(M8_UM8_0_GP34_0_GenProp8_15_line2, M8_UM8_0_GP34_0_GenProp8_15_line3, M8_PropYbus_7);
and2 M8_UM8_0_GP34_1_GenProp8_0(YAbus_8, YBbus_8, M8_GenYbus_8);
and2 M8_UM8_0_GP34_1_GenProp8_1(YAbus_9, YBbus_9, M8_GenYbus_9);
and2 M8_UM8_0_GP34_1_GenProp8_2(YAbus_10, YBbus_10, M8_GenYbus_10);
and2 M8_UM8_0_GP34_1_GenProp8_3(YAbus_11, YBbus_11, M8_GenYbus_11);
and2 M8_UM8_0_GP34_1_GenProp8_4(YAbus_12, YBbus_12, M8_GenYbus_12);
and2 M8_UM8_0_GP34_1_GenProp8_5(YAbus_13, YBbus_13, M8_GenYbus_13);
and2 M8_UM8_0_GP34_1_GenProp8_6(YAbus_14, YBbus_14, M8_GenYbus_14);
and2 M8_UM8_0_GP34_1_GenProp8_7(YAbus_15, YBbus_15, M8_GenYbus_15);
inv M8_UM8_0_GP34_1_GenProp8_8_Xo0(YAbus_8, M8_UM8_0_GP34_1_GenProp8_8_NotA);
inv M8_UM8_0_GP34_1_GenProp8_8_Xo1(YBbus_8, M8_UM8_0_GP34_1_GenProp8_8_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_8_Xo2(M8_UM8_0_GP34_1_GenProp8_8_NotA, YBbus_8, M8_UM8_0_GP34_1_GenProp8_8_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_8_Xo3(M8_UM8_0_GP34_1_GenProp8_8_NotB, YAbus_8, M8_UM8_0_GP34_1_GenProp8_8_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_8_Xo4(M8_UM8_0_GP34_1_GenProp8_8_line2, M8_UM8_0_GP34_1_GenProp8_8_line3, M8_PropYbus_8);
inv M8_UM8_0_GP34_1_GenProp8_9_Xo0(YAbus_9, M8_UM8_0_GP34_1_GenProp8_9_NotA);
inv M8_UM8_0_GP34_1_GenProp8_9_Xo1(YBbus_9, M8_UM8_0_GP34_1_GenProp8_9_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_9_Xo2(M8_UM8_0_GP34_1_GenProp8_9_NotA, YBbus_9, M8_UM8_0_GP34_1_GenProp8_9_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_9_Xo3(M8_UM8_0_GP34_1_GenProp8_9_NotB, YAbus_9, M8_UM8_0_GP34_1_GenProp8_9_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_9_Xo4(M8_UM8_0_GP34_1_GenProp8_9_line2, M8_UM8_0_GP34_1_GenProp8_9_line3, M8_PropYbus_9);
inv M8_UM8_0_GP34_1_GenProp8_10_Xo0(YAbus_10, M8_UM8_0_GP34_1_GenProp8_10_NotA);
inv M8_UM8_0_GP34_1_GenProp8_10_Xo1(YBbus_10, M8_UM8_0_GP34_1_GenProp8_10_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_10_Xo2(M8_UM8_0_GP34_1_GenProp8_10_NotA, YBbus_10, M8_UM8_0_GP34_1_GenProp8_10_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_10_Xo3(M8_UM8_0_GP34_1_GenProp8_10_NotB, YAbus_10, M8_UM8_0_GP34_1_GenProp8_10_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_10_Xo4(M8_UM8_0_GP34_1_GenProp8_10_line2, M8_UM8_0_GP34_1_GenProp8_10_line3, M8_PropYbus_10);
inv M8_UM8_0_GP34_1_GenProp8_11_Xo0(YAbus_11, M8_UM8_0_GP34_1_GenProp8_11_NotA);
inv M8_UM8_0_GP34_1_GenProp8_11_Xo1(YBbus_11, M8_UM8_0_GP34_1_GenProp8_11_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_11_Xo2(M8_UM8_0_GP34_1_GenProp8_11_NotA, YBbus_11, M8_UM8_0_GP34_1_GenProp8_11_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_11_Xo3(M8_UM8_0_GP34_1_GenProp8_11_NotB, YAbus_11, M8_UM8_0_GP34_1_GenProp8_11_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_11_Xo4(M8_UM8_0_GP34_1_GenProp8_11_line2, M8_UM8_0_GP34_1_GenProp8_11_line3, M8_PropYbus_11);
inv M8_UM8_0_GP34_1_GenProp8_12_Xo0(YAbus_12, M8_UM8_0_GP34_1_GenProp8_12_NotA);
inv M8_UM8_0_GP34_1_GenProp8_12_Xo1(YBbus_12, M8_UM8_0_GP34_1_GenProp8_12_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_12_Xo2(M8_UM8_0_GP34_1_GenProp8_12_NotA, YBbus_12, M8_UM8_0_GP34_1_GenProp8_12_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_12_Xo3(M8_UM8_0_GP34_1_GenProp8_12_NotB, YAbus_12, M8_UM8_0_GP34_1_GenProp8_12_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_12_Xo4(M8_UM8_0_GP34_1_GenProp8_12_line2, M8_UM8_0_GP34_1_GenProp8_12_line3, M8_PropYbus_12);
inv M8_UM8_0_GP34_1_GenProp8_13_Xo0(YAbus_13, M8_UM8_0_GP34_1_GenProp8_13_NotA);
inv M8_UM8_0_GP34_1_GenProp8_13_Xo1(YBbus_13, M8_UM8_0_GP34_1_GenProp8_13_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_13_Xo2(M8_UM8_0_GP34_1_GenProp8_13_NotA, YBbus_13, M8_UM8_0_GP34_1_GenProp8_13_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_13_Xo3(M8_UM8_0_GP34_1_GenProp8_13_NotB, YAbus_13, M8_UM8_0_GP34_1_GenProp8_13_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_13_Xo4(M8_UM8_0_GP34_1_GenProp8_13_line2, M8_UM8_0_GP34_1_GenProp8_13_line3, M8_PropYbus_13);
inv M8_UM8_0_GP34_1_GenProp8_14_Xo0(YAbus_14, M8_UM8_0_GP34_1_GenProp8_14_NotA);
inv M8_UM8_0_GP34_1_GenProp8_14_Xo1(YBbus_14, M8_UM8_0_GP34_1_GenProp8_14_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_14_Xo2(M8_UM8_0_GP34_1_GenProp8_14_NotA, YBbus_14, M8_UM8_0_GP34_1_GenProp8_14_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_14_Xo3(M8_UM8_0_GP34_1_GenProp8_14_NotB, YAbus_14, M8_UM8_0_GP34_1_GenProp8_14_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_14_Xo4(M8_UM8_0_GP34_1_GenProp8_14_line2, M8_UM8_0_GP34_1_GenProp8_14_line3, M8_PropYbus_14);
inv M8_UM8_0_GP34_1_GenProp8_15_Xo0(YAbus_15, M8_UM8_0_GP34_1_GenProp8_15_NotA);
inv M8_UM8_0_GP34_1_GenProp8_15_Xo1(YBbus_15, M8_UM8_0_GP34_1_GenProp8_15_NotB);
nand2 M8_UM8_0_GP34_1_GenProp8_15_Xo2(M8_UM8_0_GP34_1_GenProp8_15_NotA, YBbus_15, M8_UM8_0_GP34_1_GenProp8_15_line2);
nand2 M8_UM8_0_GP34_1_GenProp8_15_Xo3(M8_UM8_0_GP34_1_GenProp8_15_NotB, YAbus_15, M8_UM8_0_GP34_1_GenProp8_15_line3);
nand2 M8_UM8_0_GP34_1_GenProp8_15_Xo4(M8_UM8_0_GP34_1_GenProp8_15_line2, M8_UM8_0_GP34_1_GenProp8_15_line3, M8_PropYbus_15);
and2 M8_UM8_0_GP34_2_GenProp8_0(YAbus_16, YBbus_16, M8_GenYbus_16);
and2 M8_UM8_0_GP34_2_GenProp8_1(YAbus_17, YBbus_17, M8_GenYbus_17);
and2 M8_UM8_0_GP34_2_GenProp8_2(YAbus_18, YBbus_18, M8_GenYbus_18);
and2 M8_UM8_0_GP34_2_GenProp8_3(YAbus_19, YBbus_19, M8_GenYbus_19);
and2 M8_UM8_0_GP34_2_GenProp8_4(YAbus_20, YBbus_20, M8_GenYbus_20);
and2 M8_UM8_0_GP34_2_GenProp8_5(YAbus_21, YBbus_21, M8_GenYbus_21);
and2 M8_UM8_0_GP34_2_GenProp8_6(YAbus_22, YBbus_22, M8_GenYbus_22);
and2 M8_UM8_0_GP34_2_GenProp8_7(YAbus_23, YBbus_23, M8_GenYbus_23);
inv M8_UM8_0_GP34_2_GenProp8_8_Xo0(YAbus_16, M8_UM8_0_GP34_2_GenProp8_8_NotA);
inv M8_UM8_0_GP34_2_GenProp8_8_Xo1(YBbus_16, M8_UM8_0_GP34_2_GenProp8_8_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_8_Xo2(M8_UM8_0_GP34_2_GenProp8_8_NotA, YBbus_16, M8_UM8_0_GP34_2_GenProp8_8_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_8_Xo3(M8_UM8_0_GP34_2_GenProp8_8_NotB, YAbus_16, M8_UM8_0_GP34_2_GenProp8_8_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_8_Xo4(M8_UM8_0_GP34_2_GenProp8_8_line2, M8_UM8_0_GP34_2_GenProp8_8_line3, M8_PropYbus_16);
inv M8_UM8_0_GP34_2_GenProp8_9_Xo0(YAbus_17, M8_UM8_0_GP34_2_GenProp8_9_NotA);
inv M8_UM8_0_GP34_2_GenProp8_9_Xo1(YBbus_17, M8_UM8_0_GP34_2_GenProp8_9_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_9_Xo2(M8_UM8_0_GP34_2_GenProp8_9_NotA, YBbus_17, M8_UM8_0_GP34_2_GenProp8_9_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_9_Xo3(M8_UM8_0_GP34_2_GenProp8_9_NotB, YAbus_17, M8_UM8_0_GP34_2_GenProp8_9_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_9_Xo4(M8_UM8_0_GP34_2_GenProp8_9_line2, M8_UM8_0_GP34_2_GenProp8_9_line3, M8_PropYbus_17);
inv M8_UM8_0_GP34_2_GenProp8_10_Xo0(YAbus_18, M8_UM8_0_GP34_2_GenProp8_10_NotA);
inv M8_UM8_0_GP34_2_GenProp8_10_Xo1(YBbus_18, M8_UM8_0_GP34_2_GenProp8_10_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_10_Xo2(M8_UM8_0_GP34_2_GenProp8_10_NotA, YBbus_18, M8_UM8_0_GP34_2_GenProp8_10_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_10_Xo3(M8_UM8_0_GP34_2_GenProp8_10_NotB, YAbus_18, M8_UM8_0_GP34_2_GenProp8_10_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_10_Xo4(M8_UM8_0_GP34_2_GenProp8_10_line2, M8_UM8_0_GP34_2_GenProp8_10_line3, M8_PropYbus_18);
inv M8_UM8_0_GP34_2_GenProp8_11_Xo0(YAbus_19, M8_UM8_0_GP34_2_GenProp8_11_NotA);
inv M8_UM8_0_GP34_2_GenProp8_11_Xo1(YBbus_19, M8_UM8_0_GP34_2_GenProp8_11_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_11_Xo2(M8_UM8_0_GP34_2_GenProp8_11_NotA, YBbus_19, M8_UM8_0_GP34_2_GenProp8_11_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_11_Xo3(M8_UM8_0_GP34_2_GenProp8_11_NotB, YAbus_19, M8_UM8_0_GP34_2_GenProp8_11_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_11_Xo4(M8_UM8_0_GP34_2_GenProp8_11_line2, M8_UM8_0_GP34_2_GenProp8_11_line3, M8_PropYbus_19);
inv M8_UM8_0_GP34_2_GenProp8_12_Xo0(YAbus_20, M8_UM8_0_GP34_2_GenProp8_12_NotA);
inv M8_UM8_0_GP34_2_GenProp8_12_Xo1(YBbus_20, M8_UM8_0_GP34_2_GenProp8_12_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_12_Xo2(M8_UM8_0_GP34_2_GenProp8_12_NotA, YBbus_20, M8_UM8_0_GP34_2_GenProp8_12_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_12_Xo3(M8_UM8_0_GP34_2_GenProp8_12_NotB, YAbus_20, M8_UM8_0_GP34_2_GenProp8_12_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_12_Xo4(M8_UM8_0_GP34_2_GenProp8_12_line2, M8_UM8_0_GP34_2_GenProp8_12_line3, M8_PropYbus_20);
inv M8_UM8_0_GP34_2_GenProp8_13_Xo0(YAbus_21, M8_UM8_0_GP34_2_GenProp8_13_NotA);
inv M8_UM8_0_GP34_2_GenProp8_13_Xo1(YBbus_21, M8_UM8_0_GP34_2_GenProp8_13_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_13_Xo2(M8_UM8_0_GP34_2_GenProp8_13_NotA, YBbus_21, M8_UM8_0_GP34_2_GenProp8_13_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_13_Xo3(M8_UM8_0_GP34_2_GenProp8_13_NotB, YAbus_21, M8_UM8_0_GP34_2_GenProp8_13_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_13_Xo4(M8_UM8_0_GP34_2_GenProp8_13_line2, M8_UM8_0_GP34_2_GenProp8_13_line3, M8_PropYbus_21);
inv M8_UM8_0_GP34_2_GenProp8_14_Xo0(YAbus_22, M8_UM8_0_GP34_2_GenProp8_14_NotA);
inv M8_UM8_0_GP34_2_GenProp8_14_Xo1(YBbus_22, M8_UM8_0_GP34_2_GenProp8_14_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_14_Xo2(M8_UM8_0_GP34_2_GenProp8_14_NotA, YBbus_22, M8_UM8_0_GP34_2_GenProp8_14_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_14_Xo3(M8_UM8_0_GP34_2_GenProp8_14_NotB, YAbus_22, M8_UM8_0_GP34_2_GenProp8_14_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_14_Xo4(M8_UM8_0_GP34_2_GenProp8_14_line2, M8_UM8_0_GP34_2_GenProp8_14_line3, M8_PropYbus_22);
inv M8_UM8_0_GP34_2_GenProp8_15_Xo0(YAbus_23, M8_UM8_0_GP34_2_GenProp8_15_NotA);
inv M8_UM8_0_GP34_2_GenProp8_15_Xo1(YBbus_23, M8_UM8_0_GP34_2_GenProp8_15_NotB);
nand2 M8_UM8_0_GP34_2_GenProp8_15_Xo2(M8_UM8_0_GP34_2_GenProp8_15_NotA, YBbus_23, M8_UM8_0_GP34_2_GenProp8_15_line2);
nand2 M8_UM8_0_GP34_2_GenProp8_15_Xo3(M8_UM8_0_GP34_2_GenProp8_15_NotB, YAbus_23, M8_UM8_0_GP34_2_GenProp8_15_line3);
nand2 M8_UM8_0_GP34_2_GenProp8_15_Xo4(M8_UM8_0_GP34_2_GenProp8_15_line2, M8_UM8_0_GP34_2_GenProp8_15_line3, M8_PropYbus_23);
and2 M8_UM8_0_GP34_3_GenProp8_0(YAbus_24, YBbus_24, M8_GenYbus_24);
and2 M8_UM8_0_GP34_3_GenProp8_1(YAbus_25, YBbus_25, M8_GenYbus_25);
and2 M8_UM8_0_GP34_3_GenProp8_2(YAbus_26, YBbus_26, M8_GenYbus_26);
and2 M8_UM8_0_GP34_3_GenProp8_3(YAbus_27, YBbus_27, M8_GenYbus_27);
and2 M8_UM8_0_GP34_3_GenProp8_4(YAbus_28, YBbus_28, M8_GenYbus_28);
and2 M8_UM8_0_GP34_3_GenProp8_5(YAbus_29, YBbus_29, M8_GenYbus_29);
and2 M8_UM8_0_GP34_3_GenProp8_6(YAbus_30, YBbus_30, M8_GenYbus_30);
and2 M8_UM8_0_GP34_3_GenProp8_7(YAbus_31, YBbus_31, M8_GenYbus_31);
inv M8_UM8_0_GP34_3_GenProp8_8_Xo0(YAbus_24, M8_UM8_0_GP34_3_GenProp8_8_NotA);
inv M8_UM8_0_GP34_3_GenProp8_8_Xo1(YBbus_24, M8_UM8_0_GP34_3_GenProp8_8_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_8_Xo2(M8_UM8_0_GP34_3_GenProp8_8_NotA, YBbus_24, M8_UM8_0_GP34_3_GenProp8_8_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_8_Xo3(M8_UM8_0_GP34_3_GenProp8_8_NotB, YAbus_24, M8_UM8_0_GP34_3_GenProp8_8_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_8_Xo4(M8_UM8_0_GP34_3_GenProp8_8_line2, M8_UM8_0_GP34_3_GenProp8_8_line3, M8_PropYbus_24);
inv M8_UM8_0_GP34_3_GenProp8_9_Xo0(YAbus_25, M8_UM8_0_GP34_3_GenProp8_9_NotA);
inv M8_UM8_0_GP34_3_GenProp8_9_Xo1(YBbus_25, M8_UM8_0_GP34_3_GenProp8_9_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_9_Xo2(M8_UM8_0_GP34_3_GenProp8_9_NotA, YBbus_25, M8_UM8_0_GP34_3_GenProp8_9_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_9_Xo3(M8_UM8_0_GP34_3_GenProp8_9_NotB, YAbus_25, M8_UM8_0_GP34_3_GenProp8_9_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_9_Xo4(M8_UM8_0_GP34_3_GenProp8_9_line2, M8_UM8_0_GP34_3_GenProp8_9_line3, M8_PropYbus_25);
inv M8_UM8_0_GP34_3_GenProp8_10_Xo0(YAbus_26, M8_UM8_0_GP34_3_GenProp8_10_NotA);
inv M8_UM8_0_GP34_3_GenProp8_10_Xo1(YBbus_26, M8_UM8_0_GP34_3_GenProp8_10_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_10_Xo2(M8_UM8_0_GP34_3_GenProp8_10_NotA, YBbus_26, M8_UM8_0_GP34_3_GenProp8_10_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_10_Xo3(M8_UM8_0_GP34_3_GenProp8_10_NotB, YAbus_26, M8_UM8_0_GP34_3_GenProp8_10_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_10_Xo4(M8_UM8_0_GP34_3_GenProp8_10_line2, M8_UM8_0_GP34_3_GenProp8_10_line3, M8_PropYbus_26);
inv M8_UM8_0_GP34_3_GenProp8_11_Xo0(YAbus_27, M8_UM8_0_GP34_3_GenProp8_11_NotA);
inv M8_UM8_0_GP34_3_GenProp8_11_Xo1(YBbus_27, M8_UM8_0_GP34_3_GenProp8_11_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_11_Xo2(M8_UM8_0_GP34_3_GenProp8_11_NotA, YBbus_27, M8_UM8_0_GP34_3_GenProp8_11_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_11_Xo3(M8_UM8_0_GP34_3_GenProp8_11_NotB, YAbus_27, M8_UM8_0_GP34_3_GenProp8_11_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_11_Xo4(M8_UM8_0_GP34_3_GenProp8_11_line2, M8_UM8_0_GP34_3_GenProp8_11_line3, M8_PropYbus_27);
inv M8_UM8_0_GP34_3_GenProp8_12_Xo0(YAbus_28, M8_UM8_0_GP34_3_GenProp8_12_NotA);
inv M8_UM8_0_GP34_3_GenProp8_12_Xo1(YBbus_28, M8_UM8_0_GP34_3_GenProp8_12_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_12_Xo2(M8_UM8_0_GP34_3_GenProp8_12_NotA, YBbus_28, M8_UM8_0_GP34_3_GenProp8_12_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_12_Xo3(M8_UM8_0_GP34_3_GenProp8_12_NotB, YAbus_28, M8_UM8_0_GP34_3_GenProp8_12_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_12_Xo4(M8_UM8_0_GP34_3_GenProp8_12_line2, M8_UM8_0_GP34_3_GenProp8_12_line3, M8_PropYbus_28);
inv M8_UM8_0_GP34_3_GenProp8_13_Xo0(YAbus_29, M8_UM8_0_GP34_3_GenProp8_13_NotA);
inv M8_UM8_0_GP34_3_GenProp8_13_Xo1(YBbus_29, M8_UM8_0_GP34_3_GenProp8_13_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_13_Xo2(M8_UM8_0_GP34_3_GenProp8_13_NotA, YBbus_29, M8_UM8_0_GP34_3_GenProp8_13_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_13_Xo3(M8_UM8_0_GP34_3_GenProp8_13_NotB, YAbus_29, M8_UM8_0_GP34_3_GenProp8_13_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_13_Xo4(M8_UM8_0_GP34_3_GenProp8_13_line2, M8_UM8_0_GP34_3_GenProp8_13_line3, M8_PropYbus_29);
inv M8_UM8_0_GP34_3_GenProp8_14_Xo0(YAbus_30, M8_UM8_0_GP34_3_GenProp8_14_NotA);
inv M8_UM8_0_GP34_3_GenProp8_14_Xo1(YBbus_30, M8_UM8_0_GP34_3_GenProp8_14_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_14_Xo2(M8_UM8_0_GP34_3_GenProp8_14_NotA, YBbus_30, M8_UM8_0_GP34_3_GenProp8_14_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_14_Xo3(M8_UM8_0_GP34_3_GenProp8_14_NotB, YAbus_30, M8_UM8_0_GP34_3_GenProp8_14_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_14_Xo4(M8_UM8_0_GP34_3_GenProp8_14_line2, M8_UM8_0_GP34_3_GenProp8_14_line3, M8_PropYbus_30);
inv M8_UM8_0_GP34_3_GenProp8_15_Xo0(YAbus_31, M8_UM8_0_GP34_3_GenProp8_15_NotA);
inv M8_UM8_0_GP34_3_GenProp8_15_Xo1(YBbus_31, M8_UM8_0_GP34_3_GenProp8_15_NotB);
nand2 M8_UM8_0_GP34_3_GenProp8_15_Xo2(M8_UM8_0_GP34_3_GenProp8_15_NotA, YBbus_31, M8_UM8_0_GP34_3_GenProp8_15_line2);
nand2 M8_UM8_0_GP34_3_GenProp8_15_Xo3(M8_UM8_0_GP34_3_GenProp8_15_NotB, YAbus_31, M8_UM8_0_GP34_3_GenProp8_15_line3);
nand2 M8_UM8_0_GP34_3_GenProp8_15_Xo4(M8_UM8_0_GP34_3_GenProp8_15_line2, M8_UM8_0_GP34_3_GenProp8_15_line3, M8_PropYbus_31);
and2 M8_UM8_0_GP34_4(in38, YBbus_32, M8_GenYbus_32);
and2 M8_UM8_0_GP34_5(in38, YBbus_33, M8_GenYbus_33);
inv M8_UM8_0_GP34_6_Xo0(in38, M8_UM8_0_GP34_6_NotA);
inv M8_UM8_0_GP34_6_Xo1(YBbus_32, M8_UM8_0_GP34_6_NotB);
nand2 M8_UM8_0_GP34_6_Xo2(M8_UM8_0_GP34_6_NotA, YBbus_32, M8_UM8_0_GP34_6_line2);
nand2 M8_UM8_0_GP34_6_Xo3(M8_UM8_0_GP34_6_NotB, in38, M8_UM8_0_GP34_6_line3);
nand2 M8_UM8_0_GP34_6_Xo4(M8_UM8_0_GP34_6_line2, M8_UM8_0_GP34_6_line3, M8_PropYbus_32);
inv M8_UM8_0_GP34_7_Xo0(in38, M8_UM8_0_GP34_7_NotA);
inv M8_UM8_0_GP34_7_Xo1(YBbus_33, M8_UM8_0_GP34_7_NotB);
nand2 M8_UM8_0_GP34_7_Xo2(M8_UM8_0_GP34_7_NotA, YBbus_33, M8_UM8_0_GP34_7_line2);
nand2 M8_UM8_0_GP34_7_Xo3(M8_UM8_0_GP34_7_NotB, in38, M8_UM8_0_GP34_7_line3);
nand2 M8_UM8_0_GP34_7_Xo4(M8_UM8_0_GP34_7_line2, M8_UM8_0_GP34_7_line3, M8_PropYbus_33);
or2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_0(M8_GenYbus_0, M8_PropYbus_0, M8_dummy1_0);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_Ao2_0(M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_Ao2_1(M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_1_line0, M8_dummy0_1);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_Ao3a_0(M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_Ao3a_1(M8_PropYbus_1, M8_PropYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_Ao3a_2(M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_2_line1, M8_dummy1_1);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_Ao3a_0(M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_Ao3a_1(M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_Ao3a_2(M8_GenYbus_2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_3_line1, M8_dummy0_2);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_0(M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_1(M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_2(M8_PropYbus_2, M8_PropYbus_1, M8_PropYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_Ao4a_3(M8_GenYbus_2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_4_line2, M8_dummy1_2);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_0(M8_PropYbus_3, M8_GenYbus_2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_1(M8_PropYbus_3, M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_2(M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_Ao4a_3(M8_GenYbus_3, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_5_line2, M8_dummy0_3);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_0(M8_PropYbus_3, M8_GenYbus_2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_1(M8_PropYbus_3, M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_2(M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_3(M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_PropYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_Ao5a_4(M8_GenYbus_3, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_0_GLC4_6_line3, M8_dummy1_3);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_0(M8_PropYbus_4, M8_GenYbus_3, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_1(M8_PropYbus_4, M8_PropYbus_3, M8_GenYbus_2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line1);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_2(M8_PropYbus_4, M8_PropYbus_3, M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line2);
and5 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_3(M8_PropYbus_4, M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line3);
or5 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_Ao5a_4(M8_GenYbus_4, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_1_line3, M8_dummy0_4);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_0(M8_PropYbus_4, M8_GenYbus_3, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_1(M8_PropYbus_4, M8_PropYbus_3, M8_GenYbus_2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line1);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_2(M8_PropYbus_4, M8_PropYbus_3, M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line2);
and5 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_3(M8_PropYbus_4, M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line3);
and5 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_4(M8_PropYbus_4, M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_PropYbus_0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line4);
or6 M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_Ao6a_5(M8_GenYbus_4, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line2, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line3, M8_UM8_1_CC_0_GLC34_0_GLC9_0_GLC5_2_line4, M8_dummy1_4);
or2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_0(M8_GenYbus_5, M8_PropYbus_5, M8_dummy1_5);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_1_Ao2_0(M8_PropYbus_6, M8_GenYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_1_Ao2_1(M8_GenYbus_6, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_1_line0, M8_dummy0_6);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_Ao3a_0(M8_PropYbus_6, M8_GenYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_Ao3a_1(M8_PropYbus_6, M8_PropYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_Ao3a_2(M8_GenYbus_6, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_2_line1, M8_dummy1_6);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_Ao3a_0(M8_PropYbus_7, M8_GenYbus_6, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_Ao3a_1(M8_PropYbus_7, M8_PropYbus_6, M8_GenYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_Ao3a_2(M8_GenYbus_7, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_3_line1, M8_dummy0_7);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_0(M8_PropYbus_7, M8_GenYbus_6, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_1(M8_PropYbus_7, M8_PropYbus_6, M8_GenYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_2(M8_PropYbus_7, M8_PropYbus_6, M8_PropYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_Ao4a_3(M8_GenYbus_7, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_4_line2, M8_dummy1_7);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_0(M8_PropYbus_8, M8_GenYbus_7, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_1(M8_PropYbus_8, M8_PropYbus_7, M8_GenYbus_6, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_2(M8_PropYbus_8, M8_PropYbus_7, M8_PropYbus_6, M8_GenYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_Ao4a_3(M8_GenYbus_8, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_5_line2, M8_dummy0_8);
and2 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_0(M8_PropYbus_8, M8_GenYbus_7, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_1(M8_PropYbus_8, M8_PropYbus_7, M8_GenYbus_6, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_2(M8_PropYbus_8, M8_PropYbus_7, M8_PropYbus_6, M8_GenYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_3(M8_PropYbus_8, M8_PropYbus_7, M8_PropYbus_6, M8_PropYbus_5, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_Ao5a_4(M8_GenYbus_8, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_0_GLC9_4_GLC4_6_line3, M8_dummy1_8);
or2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_0(M8_GenYbus_9, M8_PropYbus_9, M8_dummy1_9);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_Ao2_0(M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_Ao2_1(M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_1_line0, M8_dummy0_10);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_Ao3a_0(M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_Ao3a_1(M8_PropYbus_10, M8_PropYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_Ao3a_2(M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_2_line1, M8_dummy1_10);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_Ao3a_0(M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_Ao3a_1(M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_Ao3a_2(M8_GenYbus_11, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_3_line1, M8_dummy0_11);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_0(M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_1(M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_2(M8_PropYbus_11, M8_PropYbus_10, M8_PropYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_Ao4a_3(M8_GenYbus_11, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_4_line2, M8_dummy1_11);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_0(M8_PropYbus_12, M8_GenYbus_11, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_1(M8_PropYbus_12, M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_2(M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_Ao4a_3(M8_GenYbus_12, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_5_line2, M8_dummy0_12);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_0(M8_PropYbus_12, M8_GenYbus_11, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_1(M8_PropYbus_12, M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_2(M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_3(M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_PropYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_Ao5a_4(M8_GenYbus_12, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_0_GLC4_6_line3, M8_dummy1_12);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_0(M8_PropYbus_13, M8_GenYbus_12, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_1(M8_PropYbus_13, M8_PropYbus_12, M8_GenYbus_11, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line1);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_2(M8_PropYbus_13, M8_PropYbus_12, M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line2);
and5 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_3(M8_PropYbus_13, M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line3);
or5 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_Ao5a_4(M8_GenYbus_13, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line2, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_1_line3, M8_dummy0_13);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_0(M8_PropYbus_13, M8_GenYbus_12, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_1(M8_PropYbus_13, M8_PropYbus_12, M8_GenYbus_11, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line1);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_2(M8_PropYbus_13, M8_PropYbus_12, M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line2);
and5 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_3(M8_PropYbus_13, M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line3);
and5 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_4(M8_PropYbus_13, M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_PropYbus_9, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line4);
or6 M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_Ao6a_5(M8_GenYbus_13, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line2, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line3, M8_UM8_1_CC_0_GLC34_1_GLC9_0_GLC5_2_line4, M8_dummy1_13);
or2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_0(M8_GenYbus_14, M8_PropYbus_14, M8_dummy1_14);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_1_Ao2_0(M8_PropYbus_15, M8_GenYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_1_Ao2_1(M8_GenYbus_15, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_1_line0, M8_dummy0_15);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_Ao3a_0(M8_PropYbus_15, M8_GenYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_Ao3a_1(M8_PropYbus_15, M8_PropYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_Ao3a_2(M8_GenYbus_15, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_2_line1, M8_dummy1_15);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_Ao3a_0(M8_PropYbus_16, M8_GenYbus_15, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_Ao3a_1(M8_PropYbus_16, M8_PropYbus_15, M8_GenYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_Ao3a_2(M8_GenYbus_16, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_3_line1, M8_dummy0_16);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_0(M8_PropYbus_16, M8_GenYbus_15, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_1(M8_PropYbus_16, M8_PropYbus_15, M8_GenYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_2(M8_PropYbus_16, M8_PropYbus_15, M8_PropYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_Ao4a_3(M8_GenYbus_16, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_4_line2, M8_dummy1_16);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_0(M8_PropYbus_17, M8_GenYbus_16, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_1(M8_PropYbus_17, M8_PropYbus_16, M8_GenYbus_15, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_2(M8_PropYbus_17, M8_PropYbus_16, M8_PropYbus_15, M8_GenYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_Ao4a_3(M8_GenYbus_17, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_5_line2, M8_dummy0_17);
and2 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_0(M8_PropYbus_17, M8_GenYbus_16, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_1(M8_PropYbus_17, M8_PropYbus_16, M8_GenYbus_15, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_2(M8_PropYbus_17, M8_PropYbus_16, M8_PropYbus_15, M8_GenYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_3(M8_PropYbus_17, M8_PropYbus_16, M8_PropYbus_15, M8_PropYbus_14, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_Ao5a_4(M8_GenYbus_17, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_1_GLC9_4_GLC4_6_line3, M8_dummy1_17);
or2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_0(M8_GenYbus_18, M8_PropYbus_18, M8_dummy1_18);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_Ao2_0(M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_Ao2_1(M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_1_line0, M8_dummy0_19);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_Ao3a_0(M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_Ao3a_1(M8_PropYbus_19, M8_PropYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_Ao3a_2(M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_2_line1, M8_dummy1_19);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_Ao3a_0(M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_Ao3a_1(M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_Ao3a_2(M8_GenYbus_20, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_3_line1, M8_dummy0_20);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_0(M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_1(M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_2(M8_PropYbus_20, M8_PropYbus_19, M8_PropYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_Ao4a_3(M8_GenYbus_20, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_4_line2, M8_dummy1_20);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_0(M8_PropYbus_21, M8_GenYbus_20, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_1(M8_PropYbus_21, M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_2(M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_Ao4a_3(M8_GenYbus_21, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_5_line2, M8_dummy0_21);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_0(M8_PropYbus_21, M8_GenYbus_20, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_1(M8_PropYbus_21, M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_2(M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_3(M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_PropYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_Ao5a_4(M8_GenYbus_21, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_0_GLC4_6_line3, M8_dummy1_21);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_0(M8_PropYbus_22, M8_GenYbus_21, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_1(M8_PropYbus_22, M8_PropYbus_21, M8_GenYbus_20, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line1);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_2(M8_PropYbus_22, M8_PropYbus_21, M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line2);
and5 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_3(M8_PropYbus_22, M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line3);
or5 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_Ao5a_4(M8_GenYbus_22, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line2, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_1_line3, M8_dummy0_22);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_0(M8_PropYbus_22, M8_GenYbus_21, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_1(M8_PropYbus_22, M8_PropYbus_21, M8_GenYbus_20, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line1);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_2(M8_PropYbus_22, M8_PropYbus_21, M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line2);
and5 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_3(M8_PropYbus_22, M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line3);
and5 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_4(M8_PropYbus_22, M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_PropYbus_18, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line4);
or6 M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_Ao6a_5(M8_GenYbus_22, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line2, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line3, M8_UM8_1_CC_0_GLC34_2_GLC9_0_GLC5_2_line4, M8_dummy1_22);
or2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_0(M8_GenYbus_23, M8_PropYbus_23, M8_dummy1_23);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_1_Ao2_0(M8_PropYbus_24, M8_GenYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_1_Ao2_1(M8_GenYbus_24, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_1_line0, M8_dummy0_24);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_Ao3a_0(M8_PropYbus_24, M8_GenYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_Ao3a_1(M8_PropYbus_24, M8_PropYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_Ao3a_2(M8_GenYbus_24, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_2_line1, M8_dummy1_24);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_Ao3a_0(M8_PropYbus_25, M8_GenYbus_24, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_Ao3a_1(M8_PropYbus_25, M8_PropYbus_24, M8_GenYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_Ao3a_2(M8_GenYbus_25, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_3_line1, M8_dummy0_25);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_0(M8_PropYbus_25, M8_GenYbus_24, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_1(M8_PropYbus_25, M8_PropYbus_24, M8_GenYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_2(M8_PropYbus_25, M8_PropYbus_24, M8_PropYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_Ao4a_3(M8_GenYbus_25, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_4_line2, M8_dummy1_25);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_0(M8_PropYbus_26, M8_GenYbus_25, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_1(M8_PropYbus_26, M8_PropYbus_25, M8_GenYbus_24, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_2(M8_PropYbus_26, M8_PropYbus_25, M8_PropYbus_24, M8_GenYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_Ao4a_3(M8_GenYbus_26, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_5_line2, M8_dummy0_26);
and2 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_0(M8_PropYbus_26, M8_GenYbus_25, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_1(M8_PropYbus_26, M8_PropYbus_25, M8_GenYbus_24, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_2(M8_PropYbus_26, M8_PropYbus_25, M8_PropYbus_24, M8_GenYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_3(M8_PropYbus_26, M8_PropYbus_25, M8_PropYbus_24, M8_PropYbus_23, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_Ao5a_4(M8_GenYbus_26, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_2_GLC9_4_GLC4_6_line3, M8_dummy1_26);
or2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_0(M8_GenYbus_27, M8_PropYbus_27, M8_dummy1_27);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_1_Ao2_0(M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_1_line0);
or2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_1_Ao2_1(M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_1_line0, M8_dummy0_28);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_Ao3a_0(M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line0);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_Ao3a_1(M8_PropYbus_28, M8_PropYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line1);
or3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_Ao3a_2(M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_2_line1, M8_dummy1_28);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_Ao3a_0(M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line0);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_Ao3a_1(M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line1);
or3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_Ao3a_2(M8_GenYbus_29, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_3_line1, M8_dummy0_29);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_0(M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line0);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_1(M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line1);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_2(M8_PropYbus_29, M8_PropYbus_28, M8_PropYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line2);
or4 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_Ao4a_3(M8_GenYbus_29, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line1, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_4_line2, M8_dummy1_29);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_0(M8_PropYbus_30, M8_GenYbus_29, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line0);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_1(M8_PropYbus_30, M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line1);
and4 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_2(M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line2);
or4 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_Ao4a_3(M8_GenYbus_30, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line1, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_5_line2, M8_dummy0_30);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_0(M8_PropYbus_30, M8_GenYbus_29, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line0);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_1(M8_PropYbus_30, M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line1);
and4 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_2(M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line2);
and4 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_3(M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_PropYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line3);
or5 M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_Ao5a_4(M8_GenYbus_30, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line1, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line2, M8_UM8_1_CC_0_GLC34_3_GLC5_0_GLC4_6_line3, M8_dummy1_30);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_1_Ao5a_0(M8_PropYbus_31, M8_GenYbus_30, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line0);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_1_Ao5a_1(M8_PropYbus_31, M8_PropYbus_30, M8_GenYbus_29, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line1);
and4 M8_UM8_1_CC_0_GLC34_3_GLC5_1_Ao5a_2(M8_PropYbus_31, M8_PropYbus_30, M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line2);
and5 M8_UM8_1_CC_0_GLC34_3_GLC5_1_Ao5a_3(M8_PropYbus_31, M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line3);
or5 M8_UM8_1_CC_0_GLC34_3_GLC5_1_Ao5a_4(M8_GenYbus_31, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line1, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line2, M8_UM8_1_CC_0_GLC34_3_GLC5_1_line3, M8_dummy0_31);
and2 M8_UM8_1_CC_0_GLC34_3_GLC5_2_Ao6a_0(M8_PropYbus_31, M8_GenYbus_30, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line0);
and3 M8_UM8_1_CC_0_GLC34_3_GLC5_2_Ao6a_1(M8_PropYbus_31, M8_PropYbus_30, M8_GenYbus_29, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line1);
and4 M8_UM8_1_CC_0_GLC34_3_GLC5_2_Ao6a_2(M8_PropYbus_31, M8_PropYbus_30, M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line2);
and5 M8_UM8_1_CC_0_GLC34_3_GLC5_2_Ao6a_3(M8_PropYbus_31, M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line3);
and5 M8_UM8_1_CC_0_GLC34_3_GLC5_2_Ao6a_4(M8_PropYbus_31, M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_PropYbus_27, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line4);
or6 M8_UM8_1_CC_0_GLC34_3_GLC5_2_Ao6a_5(M8_GenYbus_31, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line0, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line1, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line2, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line3, M8_UM8_1_CC_0_GLC34_3_GLC5_2_line4, M8_dummy1_31);
or2 M8_UM8_1_CC_0_GLC34_4_GLC2_0(M8_GenYbus_32, M8_PropYbus_32, M8_dummy1_32);
and2 M8_UM8_1_CC_0_GLC34_4_GLC2_1_Ao2_0(M8_PropYbus_33, M8_GenYbus_32, M8_UM8_1_CC_0_GLC34_4_GLC2_1_line0);
or2 M8_UM8_1_CC_0_GLC34_4_GLC2_1_Ao2_1(M8_GenYbus_33, M8_UM8_1_CC_0_GLC34_4_GLC2_1_line0, M8_dummy0_33);
and2 M8_UM8_1_CC_0_GLC34_4_GLC2_2_Ao3a_0(M8_PropYbus_33, M8_GenYbus_32, M8_UM8_1_CC_0_GLC34_4_GLC2_2_line0);
and2 M8_UM8_1_CC_0_GLC34_4_GLC2_2_Ao3a_1(M8_PropYbus_33, M8_PropYbus_32, M8_UM8_1_CC_0_GLC34_4_GLC2_2_line1);
or3 M8_UM8_1_CC_0_GLC34_4_GLC2_2_Ao3a_2(M8_GenYbus_33, M8_UM8_1_CC_0_GLC34_4_GLC2_2_line0, M8_UM8_1_CC_0_GLC34_4_GLC2_2_line1, M8_dummy1_33);
and5 M8_UM8_1_CC_1_CGC34_0_CBC0(M8_PropYbus_0, M8_PropYbus_1, M8_PropYbus_2, M8_PropYbus_3, M8_PropYbus_4, M8_UM8_1_CC_1_CGC34_0_Prop4_0);
and4 M8_UM8_1_CC_1_CGC34_0_CBC1(M8_PropYbus_5, M8_PropYbus_6, M8_PropYbus_7, M8_PropYbus_8, M8_UM8_1_CC_1_CGC34_0_Prop8_5);
and5 M8_UM8_1_CC_1_CGC34_0_CBC2(M8_PropYbus_9, M8_PropYbus_10, M8_PropYbus_11, M8_PropYbus_12, M8_PropYbus_13, M8_UM8_1_CC_1_CGC34_0_Prop13_9);
and4 M8_UM8_1_CC_1_CGC34_0_CBC3(M8_PropYbus_14, M8_PropYbus_15, M8_PropYbus_16, M8_PropYbus_17, M8_UM8_1_CC_1_CGC34_0_Prop17_14);
and5 M8_UM8_1_CC_1_CGC34_0_CBC4(M8_PropYbus_18, M8_PropYbus_19, M8_PropYbus_20, M8_PropYbus_21, M8_PropYbus_22, M8_UM8_1_CC_1_CGC34_0_Prop22_18);
and4 M8_UM8_1_CC_1_CGC34_0_CBC5(M8_PropYbus_23, M8_PropYbus_24, M8_PropYbus_25, M8_PropYbus_26, M8_UM8_1_CC_1_CGC34_0_Prop26_23);
and5 M8_UM8_1_CC_1_CGC34_0_CBC6(M8_PropYbus_27, M8_PropYbus_28, M8_PropYbus_29, M8_PropYbus_30, M8_PropYbus_31, M8_UM8_1_CC_1_CGC34_0_Prop31_27);
and2 M8_UM8_1_CC_1_CGC34_0_CBC7(M8_PropYbus_32, M8_PropYbus_33, M8_UM8_1_CC_1_CGC34_0_Prop33_32);
and2 M8_UM8_1_CC_1_CGC34_0_CBC8(M8_UM8_1_CC_1_CGC34_0_Prop4_0, M8_UM8_1_CC_1_CGC34_0_Prop8_5, M8_UM8_1_CC_1_CGC34_0_Prop8_0);
and2 M8_UM8_1_CC_1_CGC34_0_CBC9(M8_UM8_1_CC_1_CGC34_0_Prop13_9, M8_UM8_1_CC_1_CGC34_0_Prop17_14, M8_UM8_1_CC_1_CGC34_0_Prop17_9);
and2 M8_UM8_1_CC_1_CGC34_0_CBC10(M8_UM8_1_CC_1_CGC34_0_Prop22_18, M8_UM8_1_CC_1_CGC34_0_Prop26_23, M8_UM8_1_CC_1_CGC34_0_Prop26_18);
and2 M8_UM8_1_CC_1_CGC34_0_CBC11(M8_UM8_1_CC_1_CGC34_0_Prop31_27, M8_UM8_1_CC_1_CGC34_0_Prop33_32, M8_UM8_1_CC_1_CGC34_0_Prop33_27);
and2 M8_UM8_1_CC_1_CGC34_0_CBC12_Ao2_0(in89, M8_UM8_1_CC_1_CGC34_0_Prop4_0, M8_UM8_1_CC_1_CGC34_0_CBC12_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CBC12_Ao2_1(M8_dummy0_4, M8_UM8_1_CC_1_CGC34_0_CBC12_line0, M8_CarryOutYbus_4);
inv M8_UM8_1_CC_1_CGC34_0_CGC13_Mux0(M8_CarryOutYbus_4, M8_UM8_1_CC_1_CGC34_0_CGC13_Not_ContIn);
and2 M8_UM8_1_CC_1_CGC34_0_CGC13_Mux1(M8_dummy0_8, M8_UM8_1_CC_1_CGC34_0_CGC13_Not_ContIn, M8_UM8_1_CC_1_CGC34_0_CGC13_line1);
and2 M8_UM8_1_CC_1_CGC34_0_CGC13_Mux2(M8_dummy1_8, M8_CarryOutYbus_4, M8_UM8_1_CC_1_CGC34_0_CGC13_line2);
or2 M8_UM8_1_CC_1_CGC34_0_CGC13_Mux3(M8_UM8_1_CC_1_CGC34_0_CGC13_line1, M8_UM8_1_CC_1_CGC34_0_CGC13_line2, M8_CarryOutYbus_8);
and2 M8_UM8_1_CC_1_CGC34_0_GGC14_Ao2_0(M8_CarryOutYbus_8, M8_UM8_1_CC_1_CGC34_0_Prop13_9, M8_UM8_1_CC_1_CGC34_0_GGC14_line0);
or2 M8_UM8_1_CC_1_CGC34_0_GGC14_Ao2_1(M8_dummy0_13, M8_UM8_1_CC_1_CGC34_0_GGC14_line0, M8_CarryOutYbus_13);
and2 M8_UM8_1_CC_1_CGC34_0_CGC15_Ao2_0(M8_dummy0_13, M8_UM8_1_CC_1_CGC34_0_Prop17_14, M8_UM8_1_CC_1_CGC34_0_CGC15_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CGC15_Ao2_1(M8_dummy0_17, M8_UM8_1_CC_1_CGC34_0_CGC15_line0, M8_UM8_1_CC_1_CGC34_0_LocalCarry17_9);
and2 M8_UM8_1_CC_1_CGC34_0_CGC16_Ao2_0(M8_dummy0_4, M8_UM8_1_CC_1_CGC34_0_Prop8_5, M8_UM8_1_CC_1_CGC34_0_CGC16_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CGC16_Ao2_1(M8_dummy0_8, M8_UM8_1_CC_1_CGC34_0_CGC16_line0, M8_UM8_1_CC_1_CGC34_0_LocalCarry8_0);
and2 M8_UM8_1_CC_1_CGC34_0_CGC17_Ao3a_0(M8_UM8_1_CC_1_CGC34_0_Prop17_9, M8_UM8_1_CC_1_CGC34_0_LocalCarry8_0, M8_UM8_1_CC_1_CGC34_0_CGC17_line0);
and3 M8_UM8_1_CC_1_CGC34_0_CGC17_Ao3a_1(M8_UM8_1_CC_1_CGC34_0_Prop17_9, M8_UM8_1_CC_1_CGC34_0_Prop8_0, in89, M8_UM8_1_CC_1_CGC34_0_CGC17_line1);
or3 M8_UM8_1_CC_1_CGC34_0_CGC17_Ao3a_2(M8_UM8_1_CC_1_CGC34_0_LocalCarry17_9, M8_UM8_1_CC_1_CGC34_0_CGC17_line0, M8_UM8_1_CC_1_CGC34_0_CGC17_line1, out252);
and2 M8_UM8_1_CC_1_CGC34_0_CGC18_Ao2_0(out252, M8_UM8_1_CC_1_CGC34_0_Prop22_18, M8_UM8_1_CC_1_CGC34_0_CGC18_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CGC18_Ao2_1(M8_dummy0_22, M8_UM8_1_CC_1_CGC34_0_CGC18_line0, M8_CarryOutYbus_22);
and2 M8_UM8_1_CC_1_CGC34_0_CGC19_Ao2_0(M8_dummy0_22, M8_UM8_1_CC_1_CGC34_0_Prop26_23, M8_UM8_1_CC_1_CGC34_0_CGC19_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CGC19_Ao2_1(M8_dummy0_26, M8_UM8_1_CC_1_CGC34_0_CGC19_line0, M8_UM8_1_CC_1_CGC34_0_LocalCarry26_18);
and2 M8_UM8_1_CC_1_CGC34_0_CGC20_Ao4a_0(M8_UM8_1_CC_1_CGC34_0_Prop26_18, M8_UM8_1_CC_1_CGC34_0_LocalCarry17_9, M8_UM8_1_CC_1_CGC34_0_CGC20_line0);
and3 M8_UM8_1_CC_1_CGC34_0_CGC20_Ao4a_1(M8_UM8_1_CC_1_CGC34_0_Prop26_18, M8_UM8_1_CC_1_CGC34_0_Prop17_9, M8_UM8_1_CC_1_CGC34_0_LocalCarry8_0, M8_UM8_1_CC_1_CGC34_0_CGC20_line1);
and4 M8_UM8_1_CC_1_CGC34_0_CGC20_Ao4a_2(M8_UM8_1_CC_1_CGC34_0_Prop26_18, M8_UM8_1_CC_1_CGC34_0_Prop17_9, M8_UM8_1_CC_1_CGC34_0_Prop8_0, in89, M8_UM8_1_CC_1_CGC34_0_CGC20_line2);
or4 M8_UM8_1_CC_1_CGC34_0_CGC20_Ao4a_3(M8_UM8_1_CC_1_CGC34_0_LocalCarry26_18, M8_UM8_1_CC_1_CGC34_0_CGC20_line0, M8_UM8_1_CC_1_CGC34_0_CGC20_line1, M8_UM8_1_CC_1_CGC34_0_CGC20_line2, M8_CarryOutYbus_26);
and2 M8_UM8_1_CC_1_CGC34_0_CGC21_Ao2_0(M8_CarryOutYbus_26, M8_UM8_1_CC_1_CGC34_0_Prop31_27, M8_UM8_1_CC_1_CGC34_0_CGC21_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CGC21_Ao2_1(M8_dummy0_31, M8_UM8_1_CC_1_CGC34_0_CGC21_line0, M8_CarryOutYbus_31);
and2 M8_UM8_1_CC_1_CGC34_0_CGC22_Ao2_0(M8_dummy0_31, M8_UM8_1_CC_1_CGC34_0_Prop33_32, M8_UM8_1_CC_1_CGC34_0_CGC22_line0);
or2 M8_UM8_1_CC_1_CGC34_0_CGC22_Ao2_1(M8_dummy0_33, M8_UM8_1_CC_1_CGC34_0_CGC22_line0, M8_UM8_1_CC_1_CGC34_0_LocalCarry33_27);
and2 M8_UM8_1_CC_1_CGC34_0_CGC23_Ao5a_0(M8_UM8_1_CC_1_CGC34_0_Prop33_27, M8_UM8_1_CC_1_CGC34_0_LocalCarry26_18, M8_UM8_1_CC_1_CGC34_0_CGC23_line0);
and3 M8_UM8_1_CC_1_CGC34_0_CGC23_Ao5a_1(M8_UM8_1_CC_1_CGC34_0_Prop33_27, M8_UM8_1_CC_1_CGC34_0_Prop26_18, M8_UM8_1_CC_1_CGC34_0_LocalCarry17_9, M8_UM8_1_CC_1_CGC34_0_CGC23_line1);
and4 M8_UM8_1_CC_1_CGC34_0_CGC23_Ao5a_2(M8_UM8_1_CC_1_CGC34_0_Prop33_27, M8_UM8_1_CC_1_CGC34_0_Prop26_18, M8_UM8_1_CC_1_CGC34_0_Prop17_9, M8_UM8_1_CC_1_CGC34_0_LocalCarry8_0, M8_UM8_1_CC_1_CGC34_0_CGC23_line2);
and5 M8_UM8_1_CC_1_CGC34_0_CGC23_Ao5a_3(M8_UM8_1_CC_1_CGC34_0_Prop33_27, M8_UM8_1_CC_1_CGC34_0_Prop26_18, M8_UM8_1_CC_1_CGC34_0_Prop17_9, M8_UM8_1_CC_1_CGC34_0_Prop8_0, in89, M8_UM8_1_CC_1_CGC34_0_CGC23_line3);
or5 M8_UM8_1_CC_1_CGC34_0_CGC23_Ao5a_4(M8_UM8_1_CC_1_CGC34_0_LocalCarry33_27, M8_UM8_1_CC_1_CGC34_0_CGC23_line0, M8_UM8_1_CC_1_CGC34_0_CGC23_line1, M8_UM8_1_CC_1_CGC34_0_CGC23_line2, M8_UM8_1_CC_1_CGC34_0_CGC23_line3, M8_CarryOutYbus_33);
and2 M8_UM8_1_CC_1_CGC34_1_CB5_0_Ao2_0(M8_PropYbus_0, in89, M8_UM8_1_CC_1_CGC34_1_CB5_0_line0);
or2 M8_UM8_1_CC_1_CGC34_1_CB5_0_Ao2_1(M8_GenYbus_0, M8_UM8_1_CC_1_CGC34_1_CB5_0_line0, M8_CarryOutYbus_0);
and2 M8_UM8_1_CC_1_CGC34_1_CB5_1_Ao3a_0(M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_1_CGC34_1_CB5_1_line0);
and3 M8_UM8_1_CC_1_CGC34_1_CB5_1_Ao3a_1(M8_PropYbus_1, M8_PropYbus_0, in89, M8_UM8_1_CC_1_CGC34_1_CB5_1_line1);
or3 M8_UM8_1_CC_1_CGC34_1_CB5_1_Ao3a_2(M8_GenYbus_1, M8_UM8_1_CC_1_CGC34_1_CB5_1_line0, M8_UM8_1_CC_1_CGC34_1_CB5_1_line1, M8_CarryOutYbus_1);
and2 M8_UM8_1_CC_1_CGC34_1_CB5_2_Ao4a_0(M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_1_CGC34_1_CB5_2_line0);
and3 M8_UM8_1_CC_1_CGC34_1_CB5_2_Ao4a_1(M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_1_CGC34_1_CB5_2_line1);
and4 M8_UM8_1_CC_1_CGC34_1_CB5_2_Ao4a_2(M8_PropYbus_2, M8_PropYbus_1, M8_PropYbus_0, in89, M8_UM8_1_CC_1_CGC34_1_CB5_2_line2);
or4 M8_UM8_1_CC_1_CGC34_1_CB5_2_Ao4a_3(M8_GenYbus_2, M8_UM8_1_CC_1_CGC34_1_CB5_2_line0, M8_UM8_1_CC_1_CGC34_1_CB5_2_line1, M8_UM8_1_CC_1_CGC34_1_CB5_2_line2, M8_CarryOutYbus_2);
and2 M8_UM8_1_CC_1_CGC34_1_CB5_3_Ao5a_0(M8_PropYbus_3, M8_GenYbus_2, M8_UM8_1_CC_1_CGC34_1_CB5_3_line0);
and3 M8_UM8_1_CC_1_CGC34_1_CB5_3_Ao5a_1(M8_PropYbus_3, M8_PropYbus_2, M8_GenYbus_1, M8_UM8_1_CC_1_CGC34_1_CB5_3_line1);
and4 M8_UM8_1_CC_1_CGC34_1_CB5_3_Ao5a_2(M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_GenYbus_0, M8_UM8_1_CC_1_CGC34_1_CB5_3_line2);
and5 M8_UM8_1_CC_1_CGC34_1_CB5_3_Ao5a_3(M8_PropYbus_3, M8_PropYbus_2, M8_PropYbus_1, M8_PropYbus_0, in89, M8_UM8_1_CC_1_CGC34_1_CB5_3_line3);
or5 M8_UM8_1_CC_1_CGC34_1_CB5_3_Ao5a_4(M8_GenYbus_3, M8_UM8_1_CC_1_CGC34_1_CB5_3_line0, M8_UM8_1_CC_1_CGC34_1_CB5_3_line1, M8_UM8_1_CC_1_CGC34_1_CB5_3_line2, M8_UM8_1_CC_1_CGC34_1_CB5_3_line3, M8_CarryOutYbus_3);
and2 M8_UM8_1_CC_1_CGC34_2_CB5_0_Ao2_0(M8_PropYbus_9, M8_CarryOutYbus_8, M8_UM8_1_CC_1_CGC34_2_CB5_0_line0);
or2 M8_UM8_1_CC_1_CGC34_2_CB5_0_Ao2_1(M8_GenYbus_9, M8_UM8_1_CC_1_CGC34_2_CB5_0_line0, M8_CarryOutYbus_9);
and2 M8_UM8_1_CC_1_CGC34_2_CB5_1_Ao3a_0(M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_1_CGC34_2_CB5_1_line0);
and3 M8_UM8_1_CC_1_CGC34_2_CB5_1_Ao3a_1(M8_PropYbus_10, M8_PropYbus_9, M8_CarryOutYbus_8, M8_UM8_1_CC_1_CGC34_2_CB5_1_line1);
or3 M8_UM8_1_CC_1_CGC34_2_CB5_1_Ao3a_2(M8_GenYbus_10, M8_UM8_1_CC_1_CGC34_2_CB5_1_line0, M8_UM8_1_CC_1_CGC34_2_CB5_1_line1, M8_CarryOutYbus_10);
and2 M8_UM8_1_CC_1_CGC34_2_CB5_2_Ao4a_0(M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_1_CGC34_2_CB5_2_line0);
and3 M8_UM8_1_CC_1_CGC34_2_CB5_2_Ao4a_1(M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_1_CGC34_2_CB5_2_line1);
and4 M8_UM8_1_CC_1_CGC34_2_CB5_2_Ao4a_2(M8_PropYbus_11, M8_PropYbus_10, M8_PropYbus_9, M8_CarryOutYbus_8, M8_UM8_1_CC_1_CGC34_2_CB5_2_line2);
or4 M8_UM8_1_CC_1_CGC34_2_CB5_2_Ao4a_3(M8_GenYbus_11, M8_UM8_1_CC_1_CGC34_2_CB5_2_line0, M8_UM8_1_CC_1_CGC34_2_CB5_2_line1, M8_UM8_1_CC_1_CGC34_2_CB5_2_line2, M8_CarryOutYbus_11);
and2 M8_UM8_1_CC_1_CGC34_2_CB5_3_Ao5a_0(M8_PropYbus_12, M8_GenYbus_11, M8_UM8_1_CC_1_CGC34_2_CB5_3_line0);
and3 M8_UM8_1_CC_1_CGC34_2_CB5_3_Ao5a_1(M8_PropYbus_12, M8_PropYbus_11, M8_GenYbus_10, M8_UM8_1_CC_1_CGC34_2_CB5_3_line1);
and4 M8_UM8_1_CC_1_CGC34_2_CB5_3_Ao5a_2(M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_GenYbus_9, M8_UM8_1_CC_1_CGC34_2_CB5_3_line2);
and5 M8_UM8_1_CC_1_CGC34_2_CB5_3_Ao5a_3(M8_PropYbus_12, M8_PropYbus_11, M8_PropYbus_10, M8_PropYbus_9, M8_CarryOutYbus_8, M8_UM8_1_CC_1_CGC34_2_CB5_3_line3);
or5 M8_UM8_1_CC_1_CGC34_2_CB5_3_Ao5a_4(M8_GenYbus_12, M8_UM8_1_CC_1_CGC34_2_CB5_3_line0, M8_UM8_1_CC_1_CGC34_2_CB5_3_line1, M8_UM8_1_CC_1_CGC34_2_CB5_3_line2, M8_UM8_1_CC_1_CGC34_2_CB5_3_line3, M8_CarryOutYbus_12);
and2 M8_UM8_1_CC_1_CGC34_3_CB5_0_Ao2_0(M8_PropYbus_18, out252, M8_UM8_1_CC_1_CGC34_3_CB5_0_line0);
or2 M8_UM8_1_CC_1_CGC34_3_CB5_0_Ao2_1(M8_GenYbus_18, M8_UM8_1_CC_1_CGC34_3_CB5_0_line0, M8_CarryOutYbus_18);
and2 M8_UM8_1_CC_1_CGC34_3_CB5_1_Ao3a_0(M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_1_CGC34_3_CB5_1_line0);
and3 M8_UM8_1_CC_1_CGC34_3_CB5_1_Ao3a_1(M8_PropYbus_19, M8_PropYbus_18, out252, M8_UM8_1_CC_1_CGC34_3_CB5_1_line1);
or3 M8_UM8_1_CC_1_CGC34_3_CB5_1_Ao3a_2(M8_GenYbus_19, M8_UM8_1_CC_1_CGC34_3_CB5_1_line0, M8_UM8_1_CC_1_CGC34_3_CB5_1_line1, M8_CarryOutYbus_19);
and2 M8_UM8_1_CC_1_CGC34_3_CB5_2_Ao4a_0(M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_1_CGC34_3_CB5_2_line0);
and3 M8_UM8_1_CC_1_CGC34_3_CB5_2_Ao4a_1(M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_1_CGC34_3_CB5_2_line1);
and4 M8_UM8_1_CC_1_CGC34_3_CB5_2_Ao4a_2(M8_PropYbus_20, M8_PropYbus_19, M8_PropYbus_18, out252, M8_UM8_1_CC_1_CGC34_3_CB5_2_line2);
or4 M8_UM8_1_CC_1_CGC34_3_CB5_2_Ao4a_3(M8_GenYbus_20, M8_UM8_1_CC_1_CGC34_3_CB5_2_line0, M8_UM8_1_CC_1_CGC34_3_CB5_2_line1, M8_UM8_1_CC_1_CGC34_3_CB5_2_line2, M8_CarryOutYbus_20);
and2 M8_UM8_1_CC_1_CGC34_3_CB5_3_Ao5a_0(M8_PropYbus_21, M8_GenYbus_20, M8_UM8_1_CC_1_CGC34_3_CB5_3_line0);
and3 M8_UM8_1_CC_1_CGC34_3_CB5_3_Ao5a_1(M8_PropYbus_21, M8_PropYbus_20, M8_GenYbus_19, M8_UM8_1_CC_1_CGC34_3_CB5_3_line1);
and4 M8_UM8_1_CC_1_CGC34_3_CB5_3_Ao5a_2(M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_GenYbus_18, M8_UM8_1_CC_1_CGC34_3_CB5_3_line2);
and5 M8_UM8_1_CC_1_CGC34_3_CB5_3_Ao5a_3(M8_PropYbus_21, M8_PropYbus_20, M8_PropYbus_19, M8_PropYbus_18, out252, M8_UM8_1_CC_1_CGC34_3_CB5_3_line3);
or5 M8_UM8_1_CC_1_CGC34_3_CB5_3_Ao5a_4(M8_GenYbus_21, M8_UM8_1_CC_1_CGC34_3_CB5_3_line0, M8_UM8_1_CC_1_CGC34_3_CB5_3_line1, M8_UM8_1_CC_1_CGC34_3_CB5_3_line2, M8_UM8_1_CC_1_CGC34_3_CB5_3_line3, M8_CarryOutYbus_21);
and2 M8_UM8_1_CC_1_CGC34_4_CB5_0_Ao2_0(M8_PropYbus_27, M8_CarryOutYbus_26, M8_UM8_1_CC_1_CGC34_4_CB5_0_line0);
or2 M8_UM8_1_CC_1_CGC34_4_CB5_0_Ao2_1(M8_GenYbus_27, M8_UM8_1_CC_1_CGC34_4_CB5_0_line0, M8_CarryOutYbus_27);
and2 M8_UM8_1_CC_1_CGC34_4_CB5_1_Ao3a_0(M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_1_CGC34_4_CB5_1_line0);
and3 M8_UM8_1_CC_1_CGC34_4_CB5_1_Ao3a_1(M8_PropYbus_28, M8_PropYbus_27, M8_CarryOutYbus_26, M8_UM8_1_CC_1_CGC34_4_CB5_1_line1);
or3 M8_UM8_1_CC_1_CGC34_4_CB5_1_Ao3a_2(M8_GenYbus_28, M8_UM8_1_CC_1_CGC34_4_CB5_1_line0, M8_UM8_1_CC_1_CGC34_4_CB5_1_line1, M8_CarryOutYbus_28);
and2 M8_UM8_1_CC_1_CGC34_4_CB5_2_Ao4a_0(M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_1_CGC34_4_CB5_2_line0);
and3 M8_UM8_1_CC_1_CGC34_4_CB5_2_Ao4a_1(M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_1_CGC34_4_CB5_2_line1);
and4 M8_UM8_1_CC_1_CGC34_4_CB5_2_Ao4a_2(M8_PropYbus_29, M8_PropYbus_28, M8_PropYbus_27, M8_CarryOutYbus_26, M8_UM8_1_CC_1_CGC34_4_CB5_2_line2);
or4 M8_UM8_1_CC_1_CGC34_4_CB5_2_Ao4a_3(M8_GenYbus_29, M8_UM8_1_CC_1_CGC34_4_CB5_2_line0, M8_UM8_1_CC_1_CGC34_4_CB5_2_line1, M8_UM8_1_CC_1_CGC34_4_CB5_2_line2, M8_CarryOutYbus_29);
and2 M8_UM8_1_CC_1_CGC34_4_CB5_3_Ao5a_0(M8_PropYbus_30, M8_GenYbus_29, M8_UM8_1_CC_1_CGC34_4_CB5_3_line0);
and3 M8_UM8_1_CC_1_CGC34_4_CB5_3_Ao5a_1(M8_PropYbus_30, M8_PropYbus_29, M8_GenYbus_28, M8_UM8_1_CC_1_CGC34_4_CB5_3_line1);
and4 M8_UM8_1_CC_1_CGC34_4_CB5_3_Ao5a_2(M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_GenYbus_27, M8_UM8_1_CC_1_CGC34_4_CB5_3_line2);
and5 M8_UM8_1_CC_1_CGC34_4_CB5_3_Ao5a_3(M8_PropYbus_30, M8_PropYbus_29, M8_PropYbus_28, M8_PropYbus_27, M8_CarryOutYbus_26, M8_UM8_1_CC_1_CGC34_4_CB5_3_line3);
or5 M8_UM8_1_CC_1_CGC34_4_CB5_3_Ao5a_4(M8_GenYbus_30, M8_UM8_1_CC_1_CGC34_4_CB5_3_line0, M8_UM8_1_CC_1_CGC34_4_CB5_3_line1, M8_UM8_1_CC_1_CGC34_4_CB5_3_line2, M8_UM8_1_CC_1_CGC34_4_CB5_3_line3, M8_CarryOutYbus_30);
inv M8_UM8_1_CC_2_Mux0(M8_CarryOutYbus_31, M8_UM8_1_CC_2_Not_ContIn);
and2 M8_UM8_1_CC_2_Mux1(M8_dummy0_33, M8_UM8_1_CC_2_Not_ContIn, M8_UM8_1_CC_2_line1);
and2 M8_UM8_1_CC_2_Mux2(M8_dummy1_33, M8_CarryOutYbus_31, M8_UM8_1_CC_2_line2);
or2 M8_UM8_1_CC_2_Mux3(M8_UM8_1_CC_2_line1, M8_UM8_1_CC_2_line2, out249);
and4 M9_UM9_0_GS0(in150, in184, in228, in240, M9_UM9_0_K0);
and4 M9_UM9_0_GS1(in210, in152, in218, in230, M9_UM9_0_K1);
and4 M9_UM9_0_GS2(in183, in182, in185, in186, M9_UM9_0_K2);
and4 M9_UM9_0_GS3(in162, in172, in188, in199, M9_UM9_0_K3);
and2 M9_UM9_0_GS4(M9_UM9_0_K0, M9_UM9_0_K1, M9_StrobeK0_1);
and2 M9_UM9_0_GS5(M9_UM9_0_K2, M9_UM9_0_K3, M9_StrobeK2_3);
inv M9_UM9_0_GS6(M9_UM9_0_K0, out404);
inv M9_UM9_0_GS7(M9_UM9_0_K1, out406);
inv M9_UM9_0_GS8(M9_UM9_0_K2, out408);
inv M9_UM9_0_GS9(M9_UM9_0_K3, out410);
inv M9_UM9_1_PCB0_Inv7_0(in3698, M9_UM9_1_Not_PCYA0bus_0);
inv M9_UM9_1_PCB0_Inv7_1(in3701, M9_UM9_1_Not_PCYA0bus_1);
inv M9_UM9_1_PCB0_Inv7_2(in4393, M9_UM9_1_Not_PCYA0bus_2);
inv M9_UM9_1_PCB0_Inv7_3(in2208, M9_UM9_1_Not_PCYA0bus_3);
inv M9_UM9_1_PCB0_Inv7_4(in1492, M9_UM9_1_Not_PCYA0bus_4);
inv M9_UM9_1_PCB0_Inv7_5(in1496, M9_UM9_1_Not_PCYA0bus_5);
inv M9_UM9_1_PCB0_Inv7_6(in1459, M9_UM9_1_Not_PCYA0bus_6);
inv M9_UM9_1_PCB1_Mux7_0_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_0_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_0_Mux1(in229, M9_UM9_1_PCB1_Mux7_0_Not_ContIn, M9_UM9_1_PCB1_Mux7_0_line1);
and2 M9_UM9_1_PCB1_Mux7_0_Mux2(in41, MuxSel, M9_UM9_1_PCB1_Mux7_0_line2);
or2 M9_UM9_1_PCB1_Mux7_0_Mux3(M9_UM9_1_PCB1_Mux7_0_line1, M9_UM9_1_PCB1_Mux7_0_line2, M9_UM9_1_PCXAtempbus_0);
inv M9_UM9_1_PCB1_Mux7_1_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_1_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_1_Mux1(in239, M9_UM9_1_PCB1_Mux7_1_Not_ContIn, M9_UM9_1_PCB1_Mux7_1_line1);
and2 M9_UM9_1_PCB1_Mux7_1_Mux2(in44, MuxSel, M9_UM9_1_PCB1_Mux7_1_line2);
or2 M9_UM9_1_PCB1_Mux7_1_Mux3(M9_UM9_1_PCB1_Mux7_1_line1, M9_UM9_1_PCB1_Mux7_1_line2, M9_UM9_1_PCXAtempbus_1);
inv M9_UM9_1_PCB1_Mux7_2_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_2_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_2_Mux1(in227, M9_UM9_1_PCB1_Mux7_2_Not_ContIn, M9_UM9_1_PCB1_Mux7_2_line1);
and2 M9_UM9_1_PCB1_Mux7_2_Mux2(in115, MuxSel, M9_UM9_1_PCB1_Mux7_2_line2);
or2 M9_UM9_1_PCB1_Mux7_2_Mux3(M9_UM9_1_PCB1_Mux7_2_line1, M9_UM9_1_PCB1_Mux7_2_line2, M9_UM9_1_PCXAtempbus_2);
inv M9_UM9_1_PCB1_Mux7_3_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_3_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_3_Mux1(in161, M9_UM9_1_PCB1_Mux7_3_Not_ContIn, M9_UM9_1_PCB1_Mux7_3_line1);
and2 M9_UM9_1_PCB1_Mux7_3_Mux2(in141, MuxSel, M9_UM9_1_PCB1_Mux7_3_line2);
or2 M9_UM9_1_PCB1_Mux7_3_Mux3(M9_UM9_1_PCB1_Mux7_3_line1, M9_UM9_1_PCB1_Mux7_3_line2, M9_UM9_1_PCXAtempbus_3);
inv M9_UM9_1_PCB1_Mux7_4_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_4_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_4_Mux1(in212, M9_UM9_1_PCB1_Mux7_4_Not_ContIn, M9_UM9_1_PCB1_Mux7_4_line1);
and2 M9_UM9_1_PCB1_Mux7_4_Mux2(vdd, MuxSel, M9_UM9_1_PCB1_Mux7_4_line2);
or2 M9_UM9_1_PCB1_Mux7_4_Mux3(M9_UM9_1_PCB1_Mux7_4_line1, M9_UM9_1_PCB1_Mux7_4_line2, M9_UM9_1_PCXAtempbus_4);
inv M9_UM9_1_PCB1_Mux7_5_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_5_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_5_Mux1(in211, M9_UM9_1_PCB1_Mux7_5_Not_ContIn, M9_UM9_1_PCB1_Mux7_5_line1);
and2 M9_UM9_1_PCB1_Mux7_5_Mux2(vdd, MuxSel, M9_UM9_1_PCB1_Mux7_5_line2);
or2 M9_UM9_1_PCB1_Mux7_5_Mux3(M9_UM9_1_PCB1_Mux7_5_line1, M9_UM9_1_PCB1_Mux7_5_line2, M9_UM9_1_PCXAtempbus_5);
inv M9_UM9_1_PCB1_Mux7_6_Mux0(MuxSel, M9_UM9_1_PCB1_Mux7_6_Not_ContIn);
and2 M9_UM9_1_PCB1_Mux7_6_Mux1(vdd, M9_UM9_1_PCB1_Mux7_6_Not_ContIn, M9_UM9_1_PCB1_Mux7_6_line1);
and2 M9_UM9_1_PCB1_Mux7_6_Mux2(vdd, MuxSel, M9_UM9_1_PCB1_Mux7_6_line2);
or2 M9_UM9_1_PCB1_Mux7_6_Mux3(M9_UM9_1_PCB1_Mux7_6_line1, M9_UM9_1_PCB1_Mux7_6_line2, M9_UM9_1_PCXAtempbus_6);
inv M9_UM9_1_PCB2_Mux7_0_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_0_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_0_Mux1(M9_UM9_1_Not_PCYA0bus_0, M9_UM9_1_PCB2_Mux7_0_Not_ContIn, M9_UM9_1_PCB2_Mux7_0_line1);
and2 M9_UM9_1_PCB2_Mux7_0_Mux2(in69, MuxSel, M9_UM9_1_PCB2_Mux7_0_line2);
or2 M9_UM9_1_PCB2_Mux7_0_Mux3(M9_UM9_1_PCB2_Mux7_0_line1, M9_UM9_1_PCB2_Mux7_0_line2, M9_PCYAbus_0);
inv M9_UM9_1_PCB2_Mux7_1_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_1_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_1_Mux1(M9_UM9_1_Not_PCYA0bus_1, M9_UM9_1_PCB2_Mux7_1_Not_ContIn, M9_UM9_1_PCB2_Mux7_1_line1);
and2 M9_UM9_1_PCB2_Mux7_1_Mux2(in70, MuxSel, M9_UM9_1_PCB2_Mux7_1_line2);
or2 M9_UM9_1_PCB2_Mux7_1_Mux3(M9_UM9_1_PCB2_Mux7_1_line1, M9_UM9_1_PCB2_Mux7_1_line2, M9_PCYAbus_1);
inv M9_UM9_1_PCB2_Mux7_2_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_2_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_2_Mux1(M9_UM9_1_Not_PCYA0bus_2, M9_UM9_1_PCB2_Mux7_2_Not_ContIn, M9_UM9_1_PCB2_Mux7_2_line1);
and2 M9_UM9_1_PCB2_Mux7_2_Mux2(in58, MuxSel, M9_UM9_1_PCB2_Mux7_2_line2);
or2 M9_UM9_1_PCB2_Mux7_2_Mux3(M9_UM9_1_PCB2_Mux7_2_line1, M9_UM9_1_PCB2_Mux7_2_line2, M9_PCYAbus_2);
inv M9_UM9_1_PCB2_Mux7_3_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_3_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_3_Mux1(M9_UM9_1_Not_PCYA0bus_3, M9_UM9_1_PCB2_Mux7_3_Not_ContIn, M9_UM9_1_PCB2_Mux7_3_line1);
and2 M9_UM9_1_PCB2_Mux7_3_Mux2(in82, MuxSel, M9_UM9_1_PCB2_Mux7_3_line2);
or2 M9_UM9_1_PCB2_Mux7_3_Mux3(M9_UM9_1_PCB2_Mux7_3_line1, M9_UM9_1_PCB2_Mux7_3_line2, M9_PCYAbus_3);
inv M9_UM9_1_PCB2_Mux7_4_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_4_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_4_Mux1(M9_UM9_1_Not_PCYA0bus_4, M9_UM9_1_PCB2_Mux7_4_Not_ContIn, M9_UM9_1_PCB2_Mux7_4_line1);
and2 M9_UM9_1_PCB2_Mux7_4_Mux2(in1455, MuxSel, M9_UM9_1_PCB2_Mux7_4_line2);
or2 M9_UM9_1_PCB2_Mux7_4_Mux3(M9_UM9_1_PCB2_Mux7_4_line1, M9_UM9_1_PCB2_Mux7_4_line2, M9_PCYAbus_4);
inv M9_UM9_1_PCB2_Mux7_5_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_5_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_5_Mux1(M9_UM9_1_Not_PCYA0bus_5, M9_UM9_1_PCB2_Mux7_5_Not_ContIn, M9_UM9_1_PCB2_Mux7_5_line1);
and2 M9_UM9_1_PCB2_Mux7_5_Mux2(in2204, MuxSel, M9_UM9_1_PCB2_Mux7_5_line2);
or2 M9_UM9_1_PCB2_Mux7_5_Mux3(M9_UM9_1_PCB2_Mux7_5_line1, M9_UM9_1_PCB2_Mux7_5_line2, M9_PCYAbus_5);
inv M9_UM9_1_PCB2_Mux7_6_Mux0(MuxSel, M9_UM9_1_PCB2_Mux7_6_Not_ContIn);
and2 M9_UM9_1_PCB2_Mux7_6_Mux1(M9_UM9_1_Not_PCYA0bus_6, M9_UM9_1_PCB2_Mux7_6_Not_ContIn, M9_UM9_1_PCB2_Mux7_6_line1);
and2 M9_UM9_1_PCB2_Mux7_6_Mux2(in114, MuxSel, M9_UM9_1_PCB2_Mux7_6_line2);
or2 M9_UM9_1_PCB2_Mux7_6_Mux3(M9_UM9_1_PCB2_Mux7_6_line1, M9_UM9_1_PCB2_Mux7_6_line2, M9_PCYAbus_6);
inv M9_UM9_1_PCB3_Mux7_0_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_0_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_0_Mux1(in198, M9_UM9_1_PCB3_Mux7_0_Not_ContIn, M9_UM9_1_PCB3_Mux7_0_line1);
and2 M9_UM9_1_PCB3_Mux7_0_Mux2(in41, MuxSel, M9_UM9_1_PCB3_Mux7_0_line2);
or2 M9_UM9_1_PCB3_Mux7_0_Mux3(M9_UM9_1_PCB3_Mux7_0_line1, M9_UM9_1_PCB3_Mux7_0_line2, M9_UM9_1_PCYBtempbus_0);
inv M9_UM9_1_PCB3_Mux7_1_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_1_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_1_Mux1(in208, M9_UM9_1_PCB3_Mux7_1_Not_ContIn, M9_UM9_1_PCB3_Mux7_1_line1);
and2 M9_UM9_1_PCB3_Mux7_1_Mux2(in44, MuxSel, M9_UM9_1_PCB3_Mux7_1_line2);
or2 M9_UM9_1_PCB3_Mux7_1_Mux3(M9_UM9_1_PCB3_Mux7_1_line1, M9_UM9_1_PCB3_Mux7_1_line2, M9_UM9_1_PCYBtempbus_1);
inv M9_UM9_1_PCB3_Mux7_2_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_2_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_2_Mux1(in197, M9_UM9_1_PCB3_Mux7_2_Not_ContIn, M9_UM9_1_PCB3_Mux7_2_line1);
and2 M9_UM9_1_PCB3_Mux7_2_Mux2(in115, MuxSel, M9_UM9_1_PCB3_Mux7_2_line2);
or2 M9_UM9_1_PCB3_Mux7_2_Mux3(M9_UM9_1_PCB3_Mux7_2_line1, M9_UM9_1_PCB3_Mux7_2_line2, M9_UM9_1_PCYBtempbus_2);
inv M9_UM9_1_PCB3_Mux7_3_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_3_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_3_Mux1(in181, M9_UM9_1_PCB3_Mux7_3_Not_ContIn, M9_UM9_1_PCB3_Mux7_3_line1);
and2 M9_UM9_1_PCB3_Mux7_3_Mux2(in141, MuxSel, M9_UM9_1_PCB3_Mux7_3_line2);
or2 M9_UM9_1_PCB3_Mux7_3_Mux3(M9_UM9_1_PCB3_Mux7_3_line1, M9_UM9_1_PCB3_Mux7_3_line2, M9_UM9_1_PCYBtempbus_3);
inv M9_UM9_1_PCB3_Mux7_4_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_4_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_4_Mux1(in165, M9_UM9_1_PCB3_Mux7_4_Not_ContIn, M9_UM9_1_PCB3_Mux7_4_line1);
and2 M9_UM9_1_PCB3_Mux7_4_Mux2(vdd, MuxSel, M9_UM9_1_PCB3_Mux7_4_line2);
or2 M9_UM9_1_PCB3_Mux7_4_Mux3(M9_UM9_1_PCB3_Mux7_4_line1, M9_UM9_1_PCB3_Mux7_4_line2, M9_UM9_1_PCYBtempbus_4);
inv M9_UM9_1_PCB3_Mux7_5_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_5_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_5_Mux1(in164, M9_UM9_1_PCB3_Mux7_5_Not_ContIn, M9_UM9_1_PCB3_Mux7_5_line1);
and2 M9_UM9_1_PCB3_Mux7_5_Mux2(vdd, MuxSel, M9_UM9_1_PCB3_Mux7_5_line2);
or2 M9_UM9_1_PCB3_Mux7_5_Mux3(M9_UM9_1_PCB3_Mux7_5_line1, M9_UM9_1_PCB3_Mux7_5_line2, M9_UM9_1_PCYBtempbus_5);
inv M9_UM9_1_PCB3_Mux7_6_Mux0(MuxSel, M9_UM9_1_PCB3_Mux7_6_Not_ContIn);
and2 M9_UM9_1_PCB3_Mux7_6_Mux1(in170, M9_UM9_1_PCB3_Mux7_6_Not_ContIn, M9_UM9_1_PCB3_Mux7_6_line1);
and2 M9_UM9_1_PCB3_Mux7_6_Mux2(vdd, MuxSel, M9_UM9_1_PCB3_Mux7_6_line2);
or2 M9_UM9_1_PCB3_Mux7_6_Mux3(M9_UM9_1_PCB3_Mux7_6_line1, M9_UM9_1_PCB3_Mux7_6_line2, M9_UM9_1_PCYBtempbus_6);
and2 M9_UM9_1_PCB4_MN0(M9_UM9_1_PCXAtempbus_4, ContBusMask, M9_PCXAbus_4);
and2 M9_UM9_1_PCB4_MN1(M9_UM9_1_PCXAtempbus_5, ContBusMask, M9_PCXAbus_5);
and2 M9_UM9_1_PCB4_MN2(M9_UM9_1_PCXAtempbus_6, ContBusMask, M9_UM9_1_PCB4_line2);
inv M9_UM9_1_PCB4_MN3(M9_UM9_1_PCB4_line2, M9_PCXAbus_6);
and2 M9_UM9_1_PCB5_MN0(M9_UM9_1_PCYBtempbus_4, ContBusMask, M9_PCYBbus_4);
and2 M9_UM9_1_PCB5_MN1(M9_UM9_1_PCYBtempbus_5, ContBusMask, M9_PCYBbus_5);
and2 M9_UM9_1_PCB5_MN2(M9_UM9_1_PCYBtempbus_6, ContBusMask, M9_UM9_1_PCB5_line2);
inv M9_UM9_1_PCB5_MN3(M9_UM9_1_PCB5_line2, M9_PCYBbus_6);
inv M9_UM9_2_ParC0_PT0_Xo0(XAbus_5, M9_UM9_2_ParC0_PT0_NotA);
inv M9_UM9_2_ParC0_PT0_Xo1(XAbus_6, M9_UM9_2_ParC0_PT0_NotB);
nand2 M9_UM9_2_ParC0_PT0_Xo2(M9_UM9_2_ParC0_PT0_NotA, XAbus_6, M9_UM9_2_ParC0_PT0_line2);
nand2 M9_UM9_2_ParC0_PT0_Xo3(M9_UM9_2_ParC0_PT0_NotB, XAbus_5, M9_UM9_2_ParC0_PT0_line3);
nand2 M9_UM9_2_ParC0_PT0_Xo4(M9_UM9_2_ParC0_PT0_line2, M9_UM9_2_ParC0_PT0_line3, M9_UM9_2_ParC0_line0);
inv M9_UM9_2_ParC0_PT1_Xo0(XAbus_7, M9_UM9_2_ParC0_PT1_NotA);
inv M9_UM9_2_ParC0_PT1_Xo1(XAbus_8, M9_UM9_2_ParC0_PT1_NotB);
nand2 M9_UM9_2_ParC0_PT1_Xo2(M9_UM9_2_ParC0_PT1_NotA, XAbus_8, M9_UM9_2_ParC0_PT1_line2);
nand2 M9_UM9_2_ParC0_PT1_Xo3(M9_UM9_2_ParC0_PT1_NotB, XAbus_7, M9_UM9_2_ParC0_PT1_line3);
nand2 M9_UM9_2_ParC0_PT1_Xo4(M9_UM9_2_ParC0_PT1_line2, M9_UM9_2_ParC0_PT1_line3, M9_UM9_2_ParC0_line1);
inv M9_UM9_2_ParC0_PT2_Xo0(XAbus_1, M9_UM9_2_ParC0_PT2_NotA);
inv M9_UM9_2_ParC0_PT2_Xo1(XAbus_2, M9_UM9_2_ParC0_PT2_NotB);
nand2 M9_UM9_2_ParC0_PT2_Xo2(M9_UM9_2_ParC0_PT2_NotA, XAbus_2, M9_UM9_2_ParC0_PT2_line2);
nand2 M9_UM9_2_ParC0_PT2_Xo3(M9_UM9_2_ParC0_PT2_NotB, XAbus_1, M9_UM9_2_ParC0_PT2_line3);
nand2 M9_UM9_2_ParC0_PT2_Xo4(M9_UM9_2_ParC0_PT2_line2, M9_UM9_2_ParC0_PT2_line3, M9_UM9_2_ParC0_line2);
inv M9_UM9_2_ParC0_PT3_Xo0(M9_UM9_1_PCXAtempbus_0, M9_UM9_2_ParC0_PT3_NotA);
inv M9_UM9_2_ParC0_PT3_Xo1(M9_UM9_1_PCXAtempbus_1, M9_UM9_2_ParC0_PT3_NotB);
nand2 M9_UM9_2_ParC0_PT3_Xo2(M9_UM9_2_ParC0_PT3_NotA, M9_UM9_1_PCXAtempbus_1, M9_UM9_2_ParC0_PT3_line2);
nand2 M9_UM9_2_ParC0_PT3_Xo3(M9_UM9_2_ParC0_PT3_NotB, M9_UM9_1_PCXAtempbus_0, M9_UM9_2_ParC0_PT3_line3);
nand2 M9_UM9_2_ParC0_PT3_Xo4(M9_UM9_2_ParC0_PT3_line2, M9_UM9_2_ParC0_PT3_line3, M9_UM9_2_ParC0_line3);
inv M9_UM9_2_ParC0_PT4_Xo0(XAbus_3, M9_UM9_2_ParC0_PT4_NotA);
inv M9_UM9_2_ParC0_PT4_Xo1(XAbus_4, M9_UM9_2_ParC0_PT4_NotB);
nand2 M9_UM9_2_ParC0_PT4_Xo2(M9_UM9_2_ParC0_PT4_NotA, XAbus_4, M9_UM9_2_ParC0_PT4_line2);
nand2 M9_UM9_2_ParC0_PT4_Xo3(M9_UM9_2_ParC0_PT4_NotB, XAbus_3, M9_UM9_2_ParC0_PT4_line3);
nand2 M9_UM9_2_ParC0_PT4_Xo4(M9_UM9_2_ParC0_PT4_line2, M9_UM9_2_ParC0_PT4_line3, M9_UM9_2_ParC0_line4);
inv M9_UM9_2_ParC0_PT5_Xo0(M9_UM9_2_ParC0_line0, M9_UM9_2_ParC0_PT5_NotA);
inv M9_UM9_2_ParC0_PT5_Xo1(M9_UM9_2_ParC0_line1, M9_UM9_2_ParC0_PT5_NotB);
nand2 M9_UM9_2_ParC0_PT5_Xo2(M9_UM9_2_ParC0_PT5_NotA, M9_UM9_2_ParC0_line1, M9_UM9_2_ParC0_PT5_line2);
nand2 M9_UM9_2_ParC0_PT5_Xo3(M9_UM9_2_ParC0_PT5_NotB, M9_UM9_2_ParC0_line0, M9_UM9_2_ParC0_PT5_line3);
nand2 M9_UM9_2_ParC0_PT5_Xo4(M9_UM9_2_ParC0_PT5_line2, M9_UM9_2_ParC0_PT5_line3, M9_UM9_2_ParC0_line5);
inv M9_UM9_2_ParC0_PT6_Xo3_0(M9_UM9_2_ParC0_line2, M9_UM9_2_ParC0_PT6_NotA);
inv M9_UM9_2_ParC0_PT6_Xo3_1(M9_UM9_2_ParC0_line3, M9_UM9_2_ParC0_PT6_NotB);
inv M9_UM9_2_ParC0_PT6_Xo3_2(M9_UM9_2_ParC0_line4, M9_UM9_2_ParC0_PT6_NotC);
and3 M9_UM9_2_ParC0_PT6_Xo3_3(M9_UM9_2_ParC0_PT6_NotA, M9_UM9_2_ParC0_PT6_NotB, M9_UM9_2_ParC0_line4, M9_UM9_2_ParC0_PT6_line3);
and3 M9_UM9_2_ParC0_PT6_Xo3_4(M9_UM9_2_ParC0_PT6_NotA, M9_UM9_2_ParC0_line3, M9_UM9_2_ParC0_PT6_NotC, M9_UM9_2_ParC0_PT6_line4);
and3 M9_UM9_2_ParC0_PT6_Xo3_5(M9_UM9_2_ParC0_line2, M9_UM9_2_ParC0_PT6_NotB, M9_UM9_2_ParC0_PT6_NotC, M9_UM9_2_ParC0_PT6_line5);
and3 M9_UM9_2_ParC0_PT6_Xo3_6(M9_UM9_2_ParC0_line2, M9_UM9_2_ParC0_line3, M9_UM9_2_ParC0_line4, M9_UM9_2_ParC0_PT6_line6);
nor2 M9_UM9_2_ParC0_PT6_Xo3_7(M9_UM9_2_ParC0_PT6_line3, M9_UM9_2_ParC0_PT6_line4, M9_UM9_2_ParC0_PT6_line7);
nor2 M9_UM9_2_ParC0_PT6_Xo3_8(M9_UM9_2_ParC0_PT6_line5, M9_UM9_2_ParC0_PT6_line6, M9_UM9_2_ParC0_PT6_line8);
nand2 M9_UM9_2_ParC0_PT6_Xo3_9(M9_UM9_2_ParC0_PT6_line7, M9_UM9_2_ParC0_PT6_line8, M9_UM9_2_ParC0_line6);
inv M9_UM9_2_ParC0_PT7_Xo0(M9_UM9_2_ParC0_line5, M9_UM9_2_ParC0_PT7_NotA);
inv M9_UM9_2_ParC0_PT7_Xo1(M9_UM9_2_ParC0_line6, M9_UM9_2_ParC0_PT7_NotB);
nand2 M9_UM9_2_ParC0_PT7_Xo2(M9_UM9_2_ParC0_PT7_NotA, M9_UM9_2_ParC0_line6, M9_UM9_2_ParC0_PT7_line2);
nand2 M9_UM9_2_ParC0_PT7_Xo3(M9_UM9_2_ParC0_PT7_NotB, M9_UM9_2_ParC0_line5, M9_UM9_2_ParC0_PT7_line3);
nand2 M9_UM9_2_ParC0_PT7_Xo4(M9_UM9_2_ParC0_PT7_line2, M9_UM9_2_ParC0_PT7_line3, M9_UM9_2_XaP0);
inv M9_UM9_2_ParC1_PT0_Xo0(XAbus_14, M9_UM9_2_ParC1_PT0_NotA);
inv M9_UM9_2_ParC1_PT0_Xo1(XAbus_15, M9_UM9_2_ParC1_PT0_NotB);
nand2 M9_UM9_2_ParC1_PT0_Xo2(M9_UM9_2_ParC1_PT0_NotA, XAbus_15, M9_UM9_2_ParC1_PT0_line2);
nand2 M9_UM9_2_ParC1_PT0_Xo3(M9_UM9_2_ParC1_PT0_NotB, XAbus_14, M9_UM9_2_ParC1_PT0_line3);
nand2 M9_UM9_2_ParC1_PT0_Xo4(M9_UM9_2_ParC1_PT0_line2, M9_UM9_2_ParC1_PT0_line3, M9_UM9_2_ParC1_line0);
inv M9_UM9_2_ParC1_PT1_Xo0(XAbus_16, M9_UM9_2_ParC1_PT1_NotA);
inv M9_UM9_2_ParC1_PT1_Xo1(XAbus_17, M9_UM9_2_ParC1_PT1_NotB);
nand2 M9_UM9_2_ParC1_PT1_Xo2(M9_UM9_2_ParC1_PT1_NotA, XAbus_17, M9_UM9_2_ParC1_PT1_line2);
nand2 M9_UM9_2_ParC1_PT1_Xo3(M9_UM9_2_ParC1_PT1_NotB, XAbus_16, M9_UM9_2_ParC1_PT1_line3);
nand2 M9_UM9_2_ParC1_PT1_Xo4(M9_UM9_2_ParC1_PT1_line2, M9_UM9_2_ParC1_PT1_line3, M9_UM9_2_ParC1_line1);
inv M9_UM9_2_ParC1_PT2_Xo0(XAbus_10, M9_UM9_2_ParC1_PT2_NotA);
inv M9_UM9_2_ParC1_PT2_Xo1(XAbus_11, M9_UM9_2_ParC1_PT2_NotB);
nand2 M9_UM9_2_ParC1_PT2_Xo2(M9_UM9_2_ParC1_PT2_NotA, XAbus_11, M9_UM9_2_ParC1_PT2_line2);
nand2 M9_UM9_2_ParC1_PT2_Xo3(M9_UM9_2_ParC1_PT2_NotB, XAbus_10, M9_UM9_2_ParC1_PT2_line3);
nand2 M9_UM9_2_ParC1_PT2_Xo4(M9_UM9_2_ParC1_PT2_line2, M9_UM9_2_ParC1_PT2_line3, M9_UM9_2_ParC1_line2);
inv M9_UM9_2_ParC1_PT3_Xo0(M9_UM9_1_PCXAtempbus_2, M9_UM9_2_ParC1_PT3_NotA);
inv M9_UM9_2_ParC1_PT3_Xo1(XAbus_9, M9_UM9_2_ParC1_PT3_NotB);
nand2 M9_UM9_2_ParC1_PT3_Xo2(M9_UM9_2_ParC1_PT3_NotA, XAbus_9, M9_UM9_2_ParC1_PT3_line2);
nand2 M9_UM9_2_ParC1_PT3_Xo3(M9_UM9_2_ParC1_PT3_NotB, M9_UM9_1_PCXAtempbus_2, M9_UM9_2_ParC1_PT3_line3);
nand2 M9_UM9_2_ParC1_PT3_Xo4(M9_UM9_2_ParC1_PT3_line2, M9_UM9_2_ParC1_PT3_line3, M9_UM9_2_ParC1_line3);
inv M9_UM9_2_ParC1_PT4_Xo0(XAbus_12, M9_UM9_2_ParC1_PT4_NotA);
inv M9_UM9_2_ParC1_PT4_Xo1(XAbus_13, M9_UM9_2_ParC1_PT4_NotB);
nand2 M9_UM9_2_ParC1_PT4_Xo2(M9_UM9_2_ParC1_PT4_NotA, XAbus_13, M9_UM9_2_ParC1_PT4_line2);
nand2 M9_UM9_2_ParC1_PT4_Xo3(M9_UM9_2_ParC1_PT4_NotB, XAbus_12, M9_UM9_2_ParC1_PT4_line3);
nand2 M9_UM9_2_ParC1_PT4_Xo4(M9_UM9_2_ParC1_PT4_line2, M9_UM9_2_ParC1_PT4_line3, M9_UM9_2_ParC1_line4);
inv M9_UM9_2_ParC1_PT5_Xo0(M9_UM9_2_ParC1_line0, M9_UM9_2_ParC1_PT5_NotA);
inv M9_UM9_2_ParC1_PT5_Xo1(M9_UM9_2_ParC1_line1, M9_UM9_2_ParC1_PT5_NotB);
nand2 M9_UM9_2_ParC1_PT5_Xo2(M9_UM9_2_ParC1_PT5_NotA, M9_UM9_2_ParC1_line1, M9_UM9_2_ParC1_PT5_line2);
nand2 M9_UM9_2_ParC1_PT5_Xo3(M9_UM9_2_ParC1_PT5_NotB, M9_UM9_2_ParC1_line0, M9_UM9_2_ParC1_PT5_line3);
nand2 M9_UM9_2_ParC1_PT5_Xo4(M9_UM9_2_ParC1_PT5_line2, M9_UM9_2_ParC1_PT5_line3, M9_UM9_2_ParC1_line5);
inv M9_UM9_2_ParC1_PT6_Xo3_0(M9_UM9_2_ParC1_line2, M9_UM9_2_ParC1_PT6_NotA);
inv M9_UM9_2_ParC1_PT6_Xo3_1(M9_UM9_2_ParC1_line3, M9_UM9_2_ParC1_PT6_NotB);
inv M9_UM9_2_ParC1_PT6_Xo3_2(M9_UM9_2_ParC1_line4, M9_UM9_2_ParC1_PT6_NotC);
and3 M9_UM9_2_ParC1_PT6_Xo3_3(M9_UM9_2_ParC1_PT6_NotA, M9_UM9_2_ParC1_PT6_NotB, M9_UM9_2_ParC1_line4, M9_UM9_2_ParC1_PT6_line3);
and3 M9_UM9_2_ParC1_PT6_Xo3_4(M9_UM9_2_ParC1_PT6_NotA, M9_UM9_2_ParC1_line3, M9_UM9_2_ParC1_PT6_NotC, M9_UM9_2_ParC1_PT6_line4);
and3 M9_UM9_2_ParC1_PT6_Xo3_5(M9_UM9_2_ParC1_line2, M9_UM9_2_ParC1_PT6_NotB, M9_UM9_2_ParC1_PT6_NotC, M9_UM9_2_ParC1_PT6_line5);
and3 M9_UM9_2_ParC1_PT6_Xo3_6(M9_UM9_2_ParC1_line2, M9_UM9_2_ParC1_line3, M9_UM9_2_ParC1_line4, M9_UM9_2_ParC1_PT6_line6);
nor2 M9_UM9_2_ParC1_PT6_Xo3_7(M9_UM9_2_ParC1_PT6_line3, M9_UM9_2_ParC1_PT6_line4, M9_UM9_2_ParC1_PT6_line7);
nor2 M9_UM9_2_ParC1_PT6_Xo3_8(M9_UM9_2_ParC1_PT6_line5, M9_UM9_2_ParC1_PT6_line6, M9_UM9_2_ParC1_PT6_line8);
nand2 M9_UM9_2_ParC1_PT6_Xo3_9(M9_UM9_2_ParC1_PT6_line7, M9_UM9_2_ParC1_PT6_line8, M9_UM9_2_ParC1_line6);
inv M9_UM9_2_ParC1_PT7_Xo0(M9_UM9_2_ParC1_line5, M9_UM9_2_ParC1_PT7_NotA);
inv M9_UM9_2_ParC1_PT7_Xo1(M9_UM9_2_ParC1_line6, M9_UM9_2_ParC1_PT7_NotB);
nand2 M9_UM9_2_ParC1_PT7_Xo2(M9_UM9_2_ParC1_PT7_NotA, M9_UM9_2_ParC1_line6, M9_UM9_2_ParC1_PT7_line2);
nand2 M9_UM9_2_ParC1_PT7_Xo3(M9_UM9_2_ParC1_PT7_NotB, M9_UM9_2_ParC1_line5, M9_UM9_2_ParC1_PT7_line3);
nand2 M9_UM9_2_ParC1_PT7_Xo4(M9_UM9_2_ParC1_PT7_line2, M9_UM9_2_ParC1_PT7_line3, M9_UM9_2_XaP1);
inv M9_UM9_2_ParC2_PT0_Xo0(XAbus_23, M9_UM9_2_ParC2_PT0_NotA);
inv M9_UM9_2_ParC2_PT0_Xo1(XAbus_24, M9_UM9_2_ParC2_PT0_NotB);
nand2 M9_UM9_2_ParC2_PT0_Xo2(M9_UM9_2_ParC2_PT0_NotA, XAbus_24, M9_UM9_2_ParC2_PT0_line2);
nand2 M9_UM9_2_ParC2_PT0_Xo3(M9_UM9_2_ParC2_PT0_NotB, XAbus_23, M9_UM9_2_ParC2_PT0_line3);
nand2 M9_UM9_2_ParC2_PT0_Xo4(M9_UM9_2_ParC2_PT0_line2, M9_UM9_2_ParC2_PT0_line3, M9_UM9_2_ParC2_line0);
inv M9_UM9_2_ParC2_PT1_Xo0(XAbus_25, M9_UM9_2_ParC2_PT1_NotA);
inv M9_UM9_2_ParC2_PT1_Xo1(XAbus_26, M9_UM9_2_ParC2_PT1_NotB);
nand2 M9_UM9_2_ParC2_PT1_Xo2(M9_UM9_2_ParC2_PT1_NotA, XAbus_26, M9_UM9_2_ParC2_PT1_line2);
nand2 M9_UM9_2_ParC2_PT1_Xo3(M9_UM9_2_ParC2_PT1_NotB, XAbus_25, M9_UM9_2_ParC2_PT1_line3);
nand2 M9_UM9_2_ParC2_PT1_Xo4(M9_UM9_2_ParC2_PT1_line2, M9_UM9_2_ParC2_PT1_line3, M9_UM9_2_ParC2_line1);
inv M9_UM9_2_ParC2_PT2_Xo0(XAbus_19, M9_UM9_2_ParC2_PT2_NotA);
inv M9_UM9_2_ParC2_PT2_Xo1(XAbus_20, M9_UM9_2_ParC2_PT2_NotB);
nand2 M9_UM9_2_ParC2_PT2_Xo2(M9_UM9_2_ParC2_PT2_NotA, XAbus_20, M9_UM9_2_ParC2_PT2_line2);
nand2 M9_UM9_2_ParC2_PT2_Xo3(M9_UM9_2_ParC2_PT2_NotB, XAbus_19, M9_UM9_2_ParC2_PT2_line3);
nand2 M9_UM9_2_ParC2_PT2_Xo4(M9_UM9_2_ParC2_PT2_line2, M9_UM9_2_ParC2_PT2_line3, M9_UM9_2_ParC2_line2);
inv M9_UM9_2_ParC2_PT3_Xo0(M9_UM9_1_PCXAtempbus_3, M9_UM9_2_ParC2_PT3_NotA);
inv M9_UM9_2_ParC2_PT3_Xo1(XAbus_18, M9_UM9_2_ParC2_PT3_NotB);
nand2 M9_UM9_2_ParC2_PT3_Xo2(M9_UM9_2_ParC2_PT3_NotA, XAbus_18, M9_UM9_2_ParC2_PT3_line2);
nand2 M9_UM9_2_ParC2_PT3_Xo3(M9_UM9_2_ParC2_PT3_NotB, M9_UM9_1_PCXAtempbus_3, M9_UM9_2_ParC2_PT3_line3);
nand2 M9_UM9_2_ParC2_PT3_Xo4(M9_UM9_2_ParC2_PT3_line2, M9_UM9_2_ParC2_PT3_line3, M9_UM9_2_ParC2_line3);
inv M9_UM9_2_ParC2_PT4_Xo0(XAbus_21, M9_UM9_2_ParC2_PT4_NotA);
inv M9_UM9_2_ParC2_PT4_Xo1(XAbus_22, M9_UM9_2_ParC2_PT4_NotB);
nand2 M9_UM9_2_ParC2_PT4_Xo2(M9_UM9_2_ParC2_PT4_NotA, XAbus_22, M9_UM9_2_ParC2_PT4_line2);
nand2 M9_UM9_2_ParC2_PT4_Xo3(M9_UM9_2_ParC2_PT4_NotB, XAbus_21, M9_UM9_2_ParC2_PT4_line3);
nand2 M9_UM9_2_ParC2_PT4_Xo4(M9_UM9_2_ParC2_PT4_line2, M9_UM9_2_ParC2_PT4_line3, M9_UM9_2_ParC2_line4);
inv M9_UM9_2_ParC2_PT5_Xo0(M9_UM9_2_ParC2_line0, M9_UM9_2_ParC2_PT5_NotA);
inv M9_UM9_2_ParC2_PT5_Xo1(M9_UM9_2_ParC2_line1, M9_UM9_2_ParC2_PT5_NotB);
nand2 M9_UM9_2_ParC2_PT5_Xo2(M9_UM9_2_ParC2_PT5_NotA, M9_UM9_2_ParC2_line1, M9_UM9_2_ParC2_PT5_line2);
nand2 M9_UM9_2_ParC2_PT5_Xo3(M9_UM9_2_ParC2_PT5_NotB, M9_UM9_2_ParC2_line0, M9_UM9_2_ParC2_PT5_line3);
nand2 M9_UM9_2_ParC2_PT5_Xo4(M9_UM9_2_ParC2_PT5_line2, M9_UM9_2_ParC2_PT5_line3, M9_UM9_2_ParC2_line5);
inv M9_UM9_2_ParC2_PT6_Xo3_0(M9_UM9_2_ParC2_line2, M9_UM9_2_ParC2_PT6_NotA);
inv M9_UM9_2_ParC2_PT6_Xo3_1(M9_UM9_2_ParC2_line3, M9_UM9_2_ParC2_PT6_NotB);
inv M9_UM9_2_ParC2_PT6_Xo3_2(M9_UM9_2_ParC2_line4, M9_UM9_2_ParC2_PT6_NotC);
and3 M9_UM9_2_ParC2_PT6_Xo3_3(M9_UM9_2_ParC2_PT6_NotA, M9_UM9_2_ParC2_PT6_NotB, M9_UM9_2_ParC2_line4, M9_UM9_2_ParC2_PT6_line3);
and3 M9_UM9_2_ParC2_PT6_Xo3_4(M9_UM9_2_ParC2_PT6_NotA, M9_UM9_2_ParC2_line3, M9_UM9_2_ParC2_PT6_NotC, M9_UM9_2_ParC2_PT6_line4);
and3 M9_UM9_2_ParC2_PT6_Xo3_5(M9_UM9_2_ParC2_line2, M9_UM9_2_ParC2_PT6_NotB, M9_UM9_2_ParC2_PT6_NotC, M9_UM9_2_ParC2_PT6_line5);
and3 M9_UM9_2_ParC2_PT6_Xo3_6(M9_UM9_2_ParC2_line2, M9_UM9_2_ParC2_line3, M9_UM9_2_ParC2_line4, M9_UM9_2_ParC2_PT6_line6);
nor2 M9_UM9_2_ParC2_PT6_Xo3_7(M9_UM9_2_ParC2_PT6_line3, M9_UM9_2_ParC2_PT6_line4, M9_UM9_2_ParC2_PT6_line7);
nor2 M9_UM9_2_ParC2_PT6_Xo3_8(M9_UM9_2_ParC2_PT6_line5, M9_UM9_2_ParC2_PT6_line6, M9_UM9_2_ParC2_PT6_line8);
nand2 M9_UM9_2_ParC2_PT6_Xo3_9(M9_UM9_2_ParC2_PT6_line7, M9_UM9_2_ParC2_PT6_line8, M9_UM9_2_ParC2_line6);
inv M9_UM9_2_ParC2_PT7_Xo0(M9_UM9_2_ParC2_line5, M9_UM9_2_ParC2_PT7_NotA);
inv M9_UM9_2_ParC2_PT7_Xo1(M9_UM9_2_ParC2_line6, M9_UM9_2_ParC2_PT7_NotB);
nand2 M9_UM9_2_ParC2_PT7_Xo2(M9_UM9_2_ParC2_PT7_NotA, M9_UM9_2_ParC2_line6, M9_UM9_2_ParC2_PT7_line2);
nand2 M9_UM9_2_ParC2_PT7_Xo3(M9_UM9_2_ParC2_PT7_NotB, M9_UM9_2_ParC2_line5, M9_UM9_2_ParC2_PT7_line3);
nand2 M9_UM9_2_ParC2_PT7_Xo4(M9_UM9_2_ParC2_PT7_line2, M9_UM9_2_ParC2_PT7_line3, M9_UM9_2_XaP2);
inv M9_UM9_2_ParC3_PT0_Xo0(M9_PCXAbus_4, M9_UM9_2_ParC3_PT0_NotA);
inv M9_UM9_2_ParC3_PT0_Xo1(M9_PCXAbus_5, M9_UM9_2_ParC3_PT0_NotB);
nand2 M9_UM9_2_ParC3_PT0_Xo2(M9_UM9_2_ParC3_PT0_NotA, M9_PCXAbus_5, M9_UM9_2_ParC3_PT0_line2);
nand2 M9_UM9_2_ParC3_PT0_Xo3(M9_UM9_2_ParC3_PT0_NotB, M9_PCXAbus_4, M9_UM9_2_ParC3_PT0_line3);
nand2 M9_UM9_2_ParC3_PT0_Xo4(M9_UM9_2_ParC3_PT0_line2, M9_UM9_2_ParC3_PT0_line3, M9_UM9_2_ParC3_line0);
inv M9_UM9_2_ParC3_PT1_Xo0(M9_PCXAbus_6, M9_UM9_2_ParC3_PT1_NotA);
inv M9_UM9_2_ParC3_PT1_Xo1(XAbus_27, M9_UM9_2_ParC3_PT1_NotB);
nand2 M9_UM9_2_ParC3_PT1_Xo2(M9_UM9_2_ParC3_PT1_NotA, XAbus_27, M9_UM9_2_ParC3_PT1_line2);
nand2 M9_UM9_2_ParC3_PT1_Xo3(M9_UM9_2_ParC3_PT1_NotB, M9_PCXAbus_6, M9_UM9_2_ParC3_PT1_line3);
nand2 M9_UM9_2_ParC3_PT1_Xo4(M9_UM9_2_ParC3_PT1_line2, M9_UM9_2_ParC3_PT1_line3, M9_UM9_2_ParC3_line1);
inv M9_UM9_2_ParC3_PT2_Xo0(XAbus_28, M9_UM9_2_ParC3_PT2_NotA);
inv M9_UM9_2_ParC3_PT2_Xo1(XAbus_29, M9_UM9_2_ParC3_PT2_NotB);
nand2 M9_UM9_2_ParC3_PT2_Xo2(M9_UM9_2_ParC3_PT2_NotA, XAbus_29, M9_UM9_2_ParC3_PT2_line2);
nand2 M9_UM9_2_ParC3_PT2_Xo3(M9_UM9_2_ParC3_PT2_NotB, XAbus_28, M9_UM9_2_ParC3_PT2_line3);
nand2 M9_UM9_2_ParC3_PT2_Xo4(M9_UM9_2_ParC3_PT2_line2, M9_UM9_2_ParC3_PT2_line3, M9_UM9_2_ParC3_line2);
inv M9_UM9_2_ParC3_PT3_Xo0(XAbus_30, M9_UM9_2_ParC3_PT3_NotA);
inv M9_UM9_2_ParC3_PT3_Xo1(XAbus_31, M9_UM9_2_ParC3_PT3_NotB);
nand2 M9_UM9_2_ParC3_PT3_Xo2(M9_UM9_2_ParC3_PT3_NotA, XAbus_31, M9_UM9_2_ParC3_PT3_line2);
nand2 M9_UM9_2_ParC3_PT3_Xo3(M9_UM9_2_ParC3_PT3_NotB, XAbus_30, M9_UM9_2_ParC3_PT3_line3);
nand2 M9_UM9_2_ParC3_PT3_Xo4(M9_UM9_2_ParC3_PT3_line2, M9_UM9_2_ParC3_PT3_line3, M9_UM9_2_ParC3_line3);
inv M9_UM9_2_ParC3_PT4_Xo3_0(M9_UM9_2_ParC3_line1, M9_UM9_2_ParC3_PT4_NotA);
inv M9_UM9_2_ParC3_PT4_Xo3_1(M9_UM9_2_ParC3_line2, M9_UM9_2_ParC3_PT4_NotB);
inv M9_UM9_2_ParC3_PT4_Xo3_2(M9_UM9_2_ParC3_line3, M9_UM9_2_ParC3_PT4_NotC);
and3 M9_UM9_2_ParC3_PT4_Xo3_3(M9_UM9_2_ParC3_PT4_NotA, M9_UM9_2_ParC3_PT4_NotB, M9_UM9_2_ParC3_line3, M9_UM9_2_ParC3_PT4_line3);
and3 M9_UM9_2_ParC3_PT4_Xo3_4(M9_UM9_2_ParC3_PT4_NotA, M9_UM9_2_ParC3_line2, M9_UM9_2_ParC3_PT4_NotC, M9_UM9_2_ParC3_PT4_line4);
and3 M9_UM9_2_ParC3_PT4_Xo3_5(M9_UM9_2_ParC3_line1, M9_UM9_2_ParC3_PT4_NotB, M9_UM9_2_ParC3_PT4_NotC, M9_UM9_2_ParC3_PT4_line5);
and3 M9_UM9_2_ParC3_PT4_Xo3_6(M9_UM9_2_ParC3_line1, M9_UM9_2_ParC3_line2, M9_UM9_2_ParC3_line3, M9_UM9_2_ParC3_PT4_line6);
nor2 M9_UM9_2_ParC3_PT4_Xo3_7(M9_UM9_2_ParC3_PT4_line3, M9_UM9_2_ParC3_PT4_line4, M9_UM9_2_ParC3_PT4_line7);
nor2 M9_UM9_2_ParC3_PT4_Xo3_8(M9_UM9_2_ParC3_PT4_line5, M9_UM9_2_ParC3_PT4_line6, M9_UM9_2_ParC3_PT4_line8);
nand2 M9_UM9_2_ParC3_PT4_Xo3_9(M9_UM9_2_ParC3_PT4_line7, M9_UM9_2_ParC3_PT4_line8, M9_UM9_2_ParC3_line4);
inv M9_UM9_2_ParC3_PT5_Xo0(M9_UM9_2_ParC3_line0, M9_UM9_2_ParC3_PT5_NotA);
inv M9_UM9_2_ParC3_PT5_Xo1(M9_UM9_2_ParC3_line4, M9_UM9_2_ParC3_PT5_NotB);
nand2 M9_UM9_2_ParC3_PT5_Xo2(M9_UM9_2_ParC3_PT5_NotA, M9_UM9_2_ParC3_line4, M9_UM9_2_ParC3_PT5_line2);
nand2 M9_UM9_2_ParC3_PT5_Xo3(M9_UM9_2_ParC3_PT5_NotB, M9_UM9_2_ParC3_line0, M9_UM9_2_ParC3_PT5_line3);
nand2 M9_UM9_2_ParC3_PT5_Xo4(M9_UM9_2_ParC3_PT5_line2, M9_UM9_2_ParC3_PT5_line3, M9_UM9_2_XaP3);
inv M9_UM9_2_ParC4_PT0_Xo0(YAbus_5, M9_UM9_2_ParC4_PT0_NotA);
inv M9_UM9_2_ParC4_PT0_Xo1(YAbus_6, M9_UM9_2_ParC4_PT0_NotB);
nand2 M9_UM9_2_ParC4_PT0_Xo2(M9_UM9_2_ParC4_PT0_NotA, YAbus_6, M9_UM9_2_ParC4_PT0_line2);
nand2 M9_UM9_2_ParC4_PT0_Xo3(M9_UM9_2_ParC4_PT0_NotB, YAbus_5, M9_UM9_2_ParC4_PT0_line3);
nand2 M9_UM9_2_ParC4_PT0_Xo4(M9_UM9_2_ParC4_PT0_line2, M9_UM9_2_ParC4_PT0_line3, M9_UM9_2_ParC4_line0);
inv M9_UM9_2_ParC4_PT1_Xo0(YAbus_7, M9_UM9_2_ParC4_PT1_NotA);
inv M9_UM9_2_ParC4_PT1_Xo1(YAbus_8, M9_UM9_2_ParC4_PT1_NotB);
nand2 M9_UM9_2_ParC4_PT1_Xo2(M9_UM9_2_ParC4_PT1_NotA, YAbus_8, M9_UM9_2_ParC4_PT1_line2);
nand2 M9_UM9_2_ParC4_PT1_Xo3(M9_UM9_2_ParC4_PT1_NotB, YAbus_7, M9_UM9_2_ParC4_PT1_line3);
nand2 M9_UM9_2_ParC4_PT1_Xo4(M9_UM9_2_ParC4_PT1_line2, M9_UM9_2_ParC4_PT1_line3, M9_UM9_2_ParC4_line1);
inv M9_UM9_2_ParC4_PT2_Xo0(YAbus_1, M9_UM9_2_ParC4_PT2_NotA);
inv M9_UM9_2_ParC4_PT2_Xo1(YAbus_2, M9_UM9_2_ParC4_PT2_NotB);
nand2 M9_UM9_2_ParC4_PT2_Xo2(M9_UM9_2_ParC4_PT2_NotA, YAbus_2, M9_UM9_2_ParC4_PT2_line2);
nand2 M9_UM9_2_ParC4_PT2_Xo3(M9_UM9_2_ParC4_PT2_NotB, YAbus_1, M9_UM9_2_ParC4_PT2_line3);
nand2 M9_UM9_2_ParC4_PT2_Xo4(M9_UM9_2_ParC4_PT2_line2, M9_UM9_2_ParC4_PT2_line3, M9_UM9_2_ParC4_line2);
inv M9_UM9_2_ParC4_PT3_Xo0(M9_PCYAbus_0, M9_UM9_2_ParC4_PT3_NotA);
inv M9_UM9_2_ParC4_PT3_Xo1(M9_PCYAbus_1, M9_UM9_2_ParC4_PT3_NotB);
nand2 M9_UM9_2_ParC4_PT3_Xo2(M9_UM9_2_ParC4_PT3_NotA, M9_PCYAbus_1, M9_UM9_2_ParC4_PT3_line2);
nand2 M9_UM9_2_ParC4_PT3_Xo3(M9_UM9_2_ParC4_PT3_NotB, M9_PCYAbus_0, M9_UM9_2_ParC4_PT3_line3);
nand2 M9_UM9_2_ParC4_PT3_Xo4(M9_UM9_2_ParC4_PT3_line2, M9_UM9_2_ParC4_PT3_line3, M9_UM9_2_ParC4_line3);
inv M9_UM9_2_ParC4_PT4_Xo0(YAbus_3, M9_UM9_2_ParC4_PT4_NotA);
inv M9_UM9_2_ParC4_PT4_Xo1(YAbus_4, M9_UM9_2_ParC4_PT4_NotB);
nand2 M9_UM9_2_ParC4_PT4_Xo2(M9_UM9_2_ParC4_PT4_NotA, YAbus_4, M9_UM9_2_ParC4_PT4_line2);
nand2 M9_UM9_2_ParC4_PT4_Xo3(M9_UM9_2_ParC4_PT4_NotB, YAbus_3, M9_UM9_2_ParC4_PT4_line3);
nand2 M9_UM9_2_ParC4_PT4_Xo4(M9_UM9_2_ParC4_PT4_line2, M9_UM9_2_ParC4_PT4_line3, M9_UM9_2_ParC4_line4);
inv M9_UM9_2_ParC4_PT5_Xo0(M9_UM9_2_ParC4_line0, M9_UM9_2_ParC4_PT5_NotA);
inv M9_UM9_2_ParC4_PT5_Xo1(M9_UM9_2_ParC4_line1, M9_UM9_2_ParC4_PT5_NotB);
nand2 M9_UM9_2_ParC4_PT5_Xo2(M9_UM9_2_ParC4_PT5_NotA, M9_UM9_2_ParC4_line1, M9_UM9_2_ParC4_PT5_line2);
nand2 M9_UM9_2_ParC4_PT5_Xo3(M9_UM9_2_ParC4_PT5_NotB, M9_UM9_2_ParC4_line0, M9_UM9_2_ParC4_PT5_line3);
nand2 M9_UM9_2_ParC4_PT5_Xo4(M9_UM9_2_ParC4_PT5_line2, M9_UM9_2_ParC4_PT5_line3, M9_UM9_2_ParC4_line5);
inv M9_UM9_2_ParC4_PT6_Xo3_0(M9_UM9_2_ParC4_line2, M9_UM9_2_ParC4_PT6_NotA);
inv M9_UM9_2_ParC4_PT6_Xo3_1(M9_UM9_2_ParC4_line3, M9_UM9_2_ParC4_PT6_NotB);
inv M9_UM9_2_ParC4_PT6_Xo3_2(M9_UM9_2_ParC4_line4, M9_UM9_2_ParC4_PT6_NotC);
and3 M9_UM9_2_ParC4_PT6_Xo3_3(M9_UM9_2_ParC4_PT6_NotA, M9_UM9_2_ParC4_PT6_NotB, M9_UM9_2_ParC4_line4, M9_UM9_2_ParC4_PT6_line3);
and3 M9_UM9_2_ParC4_PT6_Xo3_4(M9_UM9_2_ParC4_PT6_NotA, M9_UM9_2_ParC4_line3, M9_UM9_2_ParC4_PT6_NotC, M9_UM9_2_ParC4_PT6_line4);
and3 M9_UM9_2_ParC4_PT6_Xo3_5(M9_UM9_2_ParC4_line2, M9_UM9_2_ParC4_PT6_NotB, M9_UM9_2_ParC4_PT6_NotC, M9_UM9_2_ParC4_PT6_line5);
and3 M9_UM9_2_ParC4_PT6_Xo3_6(M9_UM9_2_ParC4_line2, M9_UM9_2_ParC4_line3, M9_UM9_2_ParC4_line4, M9_UM9_2_ParC4_PT6_line6);
nor2 M9_UM9_2_ParC4_PT6_Xo3_7(M9_UM9_2_ParC4_PT6_line3, M9_UM9_2_ParC4_PT6_line4, M9_UM9_2_ParC4_PT6_line7);
nor2 M9_UM9_2_ParC4_PT6_Xo3_8(M9_UM9_2_ParC4_PT6_line5, M9_UM9_2_ParC4_PT6_line6, M9_UM9_2_ParC4_PT6_line8);
nand2 M9_UM9_2_ParC4_PT6_Xo3_9(M9_UM9_2_ParC4_PT6_line7, M9_UM9_2_ParC4_PT6_line8, M9_UM9_2_ParC4_line6);
inv M9_UM9_2_ParC4_PT7_Xo0(M9_UM9_2_ParC4_line5, M9_UM9_2_ParC4_PT7_NotA);
inv M9_UM9_2_ParC4_PT7_Xo1(M9_UM9_2_ParC4_line6, M9_UM9_2_ParC4_PT7_NotB);
nand2 M9_UM9_2_ParC4_PT7_Xo2(M9_UM9_2_ParC4_PT7_NotA, M9_UM9_2_ParC4_line6, M9_UM9_2_ParC4_PT7_line2);
nand2 M9_UM9_2_ParC4_PT7_Xo3(M9_UM9_2_ParC4_PT7_NotB, M9_UM9_2_ParC4_line5, M9_UM9_2_ParC4_PT7_line3);
nand2 M9_UM9_2_ParC4_PT7_Xo4(M9_UM9_2_ParC4_PT7_line2, M9_UM9_2_ParC4_PT7_line3, M9_UM9_2_YaP0);
inv M9_UM9_2_ParC5_PT0_Xo0(YAbus_14, M9_UM9_2_ParC5_PT0_NotA);
inv M9_UM9_2_ParC5_PT0_Xo1(YAbus_15, M9_UM9_2_ParC5_PT0_NotB);
nand2 M9_UM9_2_ParC5_PT0_Xo2(M9_UM9_2_ParC5_PT0_NotA, YAbus_15, M9_UM9_2_ParC5_PT0_line2);
nand2 M9_UM9_2_ParC5_PT0_Xo3(M9_UM9_2_ParC5_PT0_NotB, YAbus_14, M9_UM9_2_ParC5_PT0_line3);
nand2 M9_UM9_2_ParC5_PT0_Xo4(M9_UM9_2_ParC5_PT0_line2, M9_UM9_2_ParC5_PT0_line3, M9_UM9_2_ParC5_line0);
inv M9_UM9_2_ParC5_PT1_Xo0(YAbus_16, M9_UM9_2_ParC5_PT1_NotA);
inv M9_UM9_2_ParC5_PT1_Xo1(YAbus_17, M9_UM9_2_ParC5_PT1_NotB);
nand2 M9_UM9_2_ParC5_PT1_Xo2(M9_UM9_2_ParC5_PT1_NotA, YAbus_17, M9_UM9_2_ParC5_PT1_line2);
nand2 M9_UM9_2_ParC5_PT1_Xo3(M9_UM9_2_ParC5_PT1_NotB, YAbus_16, M9_UM9_2_ParC5_PT1_line3);
nand2 M9_UM9_2_ParC5_PT1_Xo4(M9_UM9_2_ParC5_PT1_line2, M9_UM9_2_ParC5_PT1_line3, M9_UM9_2_ParC5_line1);
inv M9_UM9_2_ParC5_PT2_Xo0(YAbus_10, M9_UM9_2_ParC5_PT2_NotA);
inv M9_UM9_2_ParC5_PT2_Xo1(YAbus_11, M9_UM9_2_ParC5_PT2_NotB);
nand2 M9_UM9_2_ParC5_PT2_Xo2(M9_UM9_2_ParC5_PT2_NotA, YAbus_11, M9_UM9_2_ParC5_PT2_line2);
nand2 M9_UM9_2_ParC5_PT2_Xo3(M9_UM9_2_ParC5_PT2_NotB, YAbus_10, M9_UM9_2_ParC5_PT2_line3);
nand2 M9_UM9_2_ParC5_PT2_Xo4(M9_UM9_2_ParC5_PT2_line2, M9_UM9_2_ParC5_PT2_line3, M9_UM9_2_ParC5_line2);
inv M9_UM9_2_ParC5_PT3_Xo0(M9_PCYAbus_2, M9_UM9_2_ParC5_PT3_NotA);
inv M9_UM9_2_ParC5_PT3_Xo1(YAbus_9, M9_UM9_2_ParC5_PT3_NotB);
nand2 M9_UM9_2_ParC5_PT3_Xo2(M9_UM9_2_ParC5_PT3_NotA, YAbus_9, M9_UM9_2_ParC5_PT3_line2);
nand2 M9_UM9_2_ParC5_PT3_Xo3(M9_UM9_2_ParC5_PT3_NotB, M9_PCYAbus_2, M9_UM9_2_ParC5_PT3_line3);
nand2 M9_UM9_2_ParC5_PT3_Xo4(M9_UM9_2_ParC5_PT3_line2, M9_UM9_2_ParC5_PT3_line3, M9_UM9_2_ParC5_line3);
inv M9_UM9_2_ParC5_PT4_Xo0(YAbus_12, M9_UM9_2_ParC5_PT4_NotA);
inv M9_UM9_2_ParC5_PT4_Xo1(YAbus_13, M9_UM9_2_ParC5_PT4_NotB);
nand2 M9_UM9_2_ParC5_PT4_Xo2(M9_UM9_2_ParC5_PT4_NotA, YAbus_13, M9_UM9_2_ParC5_PT4_line2);
nand2 M9_UM9_2_ParC5_PT4_Xo3(M9_UM9_2_ParC5_PT4_NotB, YAbus_12, M9_UM9_2_ParC5_PT4_line3);
nand2 M9_UM9_2_ParC5_PT4_Xo4(M9_UM9_2_ParC5_PT4_line2, M9_UM9_2_ParC5_PT4_line3, M9_UM9_2_ParC5_line4);
inv M9_UM9_2_ParC5_PT5_Xo0(M9_UM9_2_ParC5_line0, M9_UM9_2_ParC5_PT5_NotA);
inv M9_UM9_2_ParC5_PT5_Xo1(M9_UM9_2_ParC5_line1, M9_UM9_2_ParC5_PT5_NotB);
nand2 M9_UM9_2_ParC5_PT5_Xo2(M9_UM9_2_ParC5_PT5_NotA, M9_UM9_2_ParC5_line1, M9_UM9_2_ParC5_PT5_line2);
nand2 M9_UM9_2_ParC5_PT5_Xo3(M9_UM9_2_ParC5_PT5_NotB, M9_UM9_2_ParC5_line0, M9_UM9_2_ParC5_PT5_line3);
nand2 M9_UM9_2_ParC5_PT5_Xo4(M9_UM9_2_ParC5_PT5_line2, M9_UM9_2_ParC5_PT5_line3, M9_UM9_2_ParC5_line5);
inv M9_UM9_2_ParC5_PT6_Xo3_0(M9_UM9_2_ParC5_line2, M9_UM9_2_ParC5_PT6_NotA);
inv M9_UM9_2_ParC5_PT6_Xo3_1(M9_UM9_2_ParC5_line3, M9_UM9_2_ParC5_PT6_NotB);
inv M9_UM9_2_ParC5_PT6_Xo3_2(M9_UM9_2_ParC5_line4, M9_UM9_2_ParC5_PT6_NotC);
and3 M9_UM9_2_ParC5_PT6_Xo3_3(M9_UM9_2_ParC5_PT6_NotA, M9_UM9_2_ParC5_PT6_NotB, M9_UM9_2_ParC5_line4, M9_UM9_2_ParC5_PT6_line3);
and3 M9_UM9_2_ParC5_PT6_Xo3_4(M9_UM9_2_ParC5_PT6_NotA, M9_UM9_2_ParC5_line3, M9_UM9_2_ParC5_PT6_NotC, M9_UM9_2_ParC5_PT6_line4);
and3 M9_UM9_2_ParC5_PT6_Xo3_5(M9_UM9_2_ParC5_line2, M9_UM9_2_ParC5_PT6_NotB, M9_UM9_2_ParC5_PT6_NotC, M9_UM9_2_ParC5_PT6_line5);
and3 M9_UM9_2_ParC5_PT6_Xo3_6(M9_UM9_2_ParC5_line2, M9_UM9_2_ParC5_line3, M9_UM9_2_ParC5_line4, M9_UM9_2_ParC5_PT6_line6);
nor2 M9_UM9_2_ParC5_PT6_Xo3_7(M9_UM9_2_ParC5_PT6_line3, M9_UM9_2_ParC5_PT6_line4, M9_UM9_2_ParC5_PT6_line7);
nor2 M9_UM9_2_ParC5_PT6_Xo3_8(M9_UM9_2_ParC5_PT6_line5, M9_UM9_2_ParC5_PT6_line6, M9_UM9_2_ParC5_PT6_line8);
nand2 M9_UM9_2_ParC5_PT6_Xo3_9(M9_UM9_2_ParC5_PT6_line7, M9_UM9_2_ParC5_PT6_line8, M9_UM9_2_ParC5_line6);
inv M9_UM9_2_ParC5_PT7_Xo0(M9_UM9_2_ParC5_line5, M9_UM9_2_ParC5_PT7_NotA);
inv M9_UM9_2_ParC5_PT7_Xo1(M9_UM9_2_ParC5_line6, M9_UM9_2_ParC5_PT7_NotB);
nand2 M9_UM9_2_ParC5_PT7_Xo2(M9_UM9_2_ParC5_PT7_NotA, M9_UM9_2_ParC5_line6, M9_UM9_2_ParC5_PT7_line2);
nand2 M9_UM9_2_ParC5_PT7_Xo3(M9_UM9_2_ParC5_PT7_NotB, M9_UM9_2_ParC5_line5, M9_UM9_2_ParC5_PT7_line3);
nand2 M9_UM9_2_ParC5_PT7_Xo4(M9_UM9_2_ParC5_PT7_line2, M9_UM9_2_ParC5_PT7_line3, M9_UM9_2_YaP1);
inv M9_UM9_2_ParC6_PT0_Xo0(YAbus_23, M9_UM9_2_ParC6_PT0_NotA);
inv M9_UM9_2_ParC6_PT0_Xo1(YAbus_24, M9_UM9_2_ParC6_PT0_NotB);
nand2 M9_UM9_2_ParC6_PT0_Xo2(M9_UM9_2_ParC6_PT0_NotA, YAbus_24, M9_UM9_2_ParC6_PT0_line2);
nand2 M9_UM9_2_ParC6_PT0_Xo3(M9_UM9_2_ParC6_PT0_NotB, YAbus_23, M9_UM9_2_ParC6_PT0_line3);
nand2 M9_UM9_2_ParC6_PT0_Xo4(M9_UM9_2_ParC6_PT0_line2, M9_UM9_2_ParC6_PT0_line3, M9_UM9_2_ParC6_line0);
inv M9_UM9_2_ParC6_PT1_Xo0(YAbus_25, M9_UM9_2_ParC6_PT1_NotA);
inv M9_UM9_2_ParC6_PT1_Xo1(YAbus_26, M9_UM9_2_ParC6_PT1_NotB);
nand2 M9_UM9_2_ParC6_PT1_Xo2(M9_UM9_2_ParC6_PT1_NotA, YAbus_26, M9_UM9_2_ParC6_PT1_line2);
nand2 M9_UM9_2_ParC6_PT1_Xo3(M9_UM9_2_ParC6_PT1_NotB, YAbus_25, M9_UM9_2_ParC6_PT1_line3);
nand2 M9_UM9_2_ParC6_PT1_Xo4(M9_UM9_2_ParC6_PT1_line2, M9_UM9_2_ParC6_PT1_line3, M9_UM9_2_ParC6_line1);
inv M9_UM9_2_ParC6_PT2_Xo0(YAbus_19, M9_UM9_2_ParC6_PT2_NotA);
inv M9_UM9_2_ParC6_PT2_Xo1(YAbus_20, M9_UM9_2_ParC6_PT2_NotB);
nand2 M9_UM9_2_ParC6_PT2_Xo2(M9_UM9_2_ParC6_PT2_NotA, YAbus_20, M9_UM9_2_ParC6_PT2_line2);
nand2 M9_UM9_2_ParC6_PT2_Xo3(M9_UM9_2_ParC6_PT2_NotB, YAbus_19, M9_UM9_2_ParC6_PT2_line3);
nand2 M9_UM9_2_ParC6_PT2_Xo4(M9_UM9_2_ParC6_PT2_line2, M9_UM9_2_ParC6_PT2_line3, M9_UM9_2_ParC6_line2);
inv M9_UM9_2_ParC6_PT3_Xo0(M9_PCYAbus_3, M9_UM9_2_ParC6_PT3_NotA);
inv M9_UM9_2_ParC6_PT3_Xo1(YAbus_18, M9_UM9_2_ParC6_PT3_NotB);
nand2 M9_UM9_2_ParC6_PT3_Xo2(M9_UM9_2_ParC6_PT3_NotA, YAbus_18, M9_UM9_2_ParC6_PT3_line2);
nand2 M9_UM9_2_ParC6_PT3_Xo3(M9_UM9_2_ParC6_PT3_NotB, M9_PCYAbus_3, M9_UM9_2_ParC6_PT3_line3);
nand2 M9_UM9_2_ParC6_PT3_Xo4(M9_UM9_2_ParC6_PT3_line2, M9_UM9_2_ParC6_PT3_line3, M9_UM9_2_ParC6_line3);
inv M9_UM9_2_ParC6_PT4_Xo0(YAbus_21, M9_UM9_2_ParC6_PT4_NotA);
inv M9_UM9_2_ParC6_PT4_Xo1(YAbus_22, M9_UM9_2_ParC6_PT4_NotB);
nand2 M9_UM9_2_ParC6_PT4_Xo2(M9_UM9_2_ParC6_PT4_NotA, YAbus_22, M9_UM9_2_ParC6_PT4_line2);
nand2 M9_UM9_2_ParC6_PT4_Xo3(M9_UM9_2_ParC6_PT4_NotB, YAbus_21, M9_UM9_2_ParC6_PT4_line3);
nand2 M9_UM9_2_ParC6_PT4_Xo4(M9_UM9_2_ParC6_PT4_line2, M9_UM9_2_ParC6_PT4_line3, M9_UM9_2_ParC6_line4);
inv M9_UM9_2_ParC6_PT5_Xo0(M9_UM9_2_ParC6_line0, M9_UM9_2_ParC6_PT5_NotA);
inv M9_UM9_2_ParC6_PT5_Xo1(M9_UM9_2_ParC6_line1, M9_UM9_2_ParC6_PT5_NotB);
nand2 M9_UM9_2_ParC6_PT5_Xo2(M9_UM9_2_ParC6_PT5_NotA, M9_UM9_2_ParC6_line1, M9_UM9_2_ParC6_PT5_line2);
nand2 M9_UM9_2_ParC6_PT5_Xo3(M9_UM9_2_ParC6_PT5_NotB, M9_UM9_2_ParC6_line0, M9_UM9_2_ParC6_PT5_line3);
nand2 M9_UM9_2_ParC6_PT5_Xo4(M9_UM9_2_ParC6_PT5_line2, M9_UM9_2_ParC6_PT5_line3, M9_UM9_2_ParC6_line5);
inv M9_UM9_2_ParC6_PT6_Xo3_0(M9_UM9_2_ParC6_line2, M9_UM9_2_ParC6_PT6_NotA);
inv M9_UM9_2_ParC6_PT6_Xo3_1(M9_UM9_2_ParC6_line3, M9_UM9_2_ParC6_PT6_NotB);
inv M9_UM9_2_ParC6_PT6_Xo3_2(M9_UM9_2_ParC6_line4, M9_UM9_2_ParC6_PT6_NotC);
and3 M9_UM9_2_ParC6_PT6_Xo3_3(M9_UM9_2_ParC6_PT6_NotA, M9_UM9_2_ParC6_PT6_NotB, M9_UM9_2_ParC6_line4, M9_UM9_2_ParC6_PT6_line3);
and3 M9_UM9_2_ParC6_PT6_Xo3_4(M9_UM9_2_ParC6_PT6_NotA, M9_UM9_2_ParC6_line3, M9_UM9_2_ParC6_PT6_NotC, M9_UM9_2_ParC6_PT6_line4);
and3 M9_UM9_2_ParC6_PT6_Xo3_5(M9_UM9_2_ParC6_line2, M9_UM9_2_ParC6_PT6_NotB, M9_UM9_2_ParC6_PT6_NotC, M9_UM9_2_ParC6_PT6_line5);
and3 M9_UM9_2_ParC6_PT6_Xo3_6(M9_UM9_2_ParC6_line2, M9_UM9_2_ParC6_line3, M9_UM9_2_ParC6_line4, M9_UM9_2_ParC6_PT6_line6);
nor2 M9_UM9_2_ParC6_PT6_Xo3_7(M9_UM9_2_ParC6_PT6_line3, M9_UM9_2_ParC6_PT6_line4, M9_UM9_2_ParC6_PT6_line7);
nor2 M9_UM9_2_ParC6_PT6_Xo3_8(M9_UM9_2_ParC6_PT6_line5, M9_UM9_2_ParC6_PT6_line6, M9_UM9_2_ParC6_PT6_line8);
nand2 M9_UM9_2_ParC6_PT6_Xo3_9(M9_UM9_2_ParC6_PT6_line7, M9_UM9_2_ParC6_PT6_line8, M9_UM9_2_ParC6_line6);
inv M9_UM9_2_ParC6_PT7_Xo0(M9_UM9_2_ParC6_line5, M9_UM9_2_ParC6_PT7_NotA);
inv M9_UM9_2_ParC6_PT7_Xo1(M9_UM9_2_ParC6_line6, M9_UM9_2_ParC6_PT7_NotB);
nand2 M9_UM9_2_ParC6_PT7_Xo2(M9_UM9_2_ParC6_PT7_NotA, M9_UM9_2_ParC6_line6, M9_UM9_2_ParC6_PT7_line2);
nand2 M9_UM9_2_ParC6_PT7_Xo3(M9_UM9_2_ParC6_PT7_NotB, M9_UM9_2_ParC6_line5, M9_UM9_2_ParC6_PT7_line3);
nand2 M9_UM9_2_ParC6_PT7_Xo4(M9_UM9_2_ParC6_PT7_line2, M9_UM9_2_ParC6_PT7_line3, M9_UM9_2_YaP2);
inv M9_UM9_2_ParC7_PT0_Xo0(M9_PCYAbus_4, M9_UM9_2_ParC7_PT0_NotA);
inv M9_UM9_2_ParC7_PT0_Xo1(M9_PCYAbus_5, M9_UM9_2_ParC7_PT0_NotB);
nand2 M9_UM9_2_ParC7_PT0_Xo2(M9_UM9_2_ParC7_PT0_NotA, M9_PCYAbus_5, M9_UM9_2_ParC7_PT0_line2);
nand2 M9_UM9_2_ParC7_PT0_Xo3(M9_UM9_2_ParC7_PT0_NotB, M9_PCYAbus_4, M9_UM9_2_ParC7_PT0_line3);
nand2 M9_UM9_2_ParC7_PT0_Xo4(M9_UM9_2_ParC7_PT0_line2, M9_UM9_2_ParC7_PT0_line3, M9_UM9_2_ParC7_line0);
inv M9_UM9_2_ParC7_PT1_Xo0(M9_PCYAbus_6, M9_UM9_2_ParC7_PT1_NotA);
inv M9_UM9_2_ParC7_PT1_Xo1(YAbus_27, M9_UM9_2_ParC7_PT1_NotB);
nand2 M9_UM9_2_ParC7_PT1_Xo2(M9_UM9_2_ParC7_PT1_NotA, YAbus_27, M9_UM9_2_ParC7_PT1_line2);
nand2 M9_UM9_2_ParC7_PT1_Xo3(M9_UM9_2_ParC7_PT1_NotB, M9_PCYAbus_6, M9_UM9_2_ParC7_PT1_line3);
nand2 M9_UM9_2_ParC7_PT1_Xo4(M9_UM9_2_ParC7_PT1_line2, M9_UM9_2_ParC7_PT1_line3, M9_UM9_2_ParC7_line1);
inv M9_UM9_2_ParC7_PT2_Xo0(YAbus_28, M9_UM9_2_ParC7_PT2_NotA);
inv M9_UM9_2_ParC7_PT2_Xo1(YAbus_29, M9_UM9_2_ParC7_PT2_NotB);
nand2 M9_UM9_2_ParC7_PT2_Xo2(M9_UM9_2_ParC7_PT2_NotA, YAbus_29, M9_UM9_2_ParC7_PT2_line2);
nand2 M9_UM9_2_ParC7_PT2_Xo3(M9_UM9_2_ParC7_PT2_NotB, YAbus_28, M9_UM9_2_ParC7_PT2_line3);
nand2 M9_UM9_2_ParC7_PT2_Xo4(M9_UM9_2_ParC7_PT2_line2, M9_UM9_2_ParC7_PT2_line3, M9_UM9_2_ParC7_line2);
inv M9_UM9_2_ParC7_PT3_Xo0(YAbus_30, M9_UM9_2_ParC7_PT3_NotA);
inv M9_UM9_2_ParC7_PT3_Xo1(YAbus_31, M9_UM9_2_ParC7_PT3_NotB);
nand2 M9_UM9_2_ParC7_PT3_Xo2(M9_UM9_2_ParC7_PT3_NotA, YAbus_31, M9_UM9_2_ParC7_PT3_line2);
nand2 M9_UM9_2_ParC7_PT3_Xo3(M9_UM9_2_ParC7_PT3_NotB, YAbus_30, M9_UM9_2_ParC7_PT3_line3);
nand2 M9_UM9_2_ParC7_PT3_Xo4(M9_UM9_2_ParC7_PT3_line2, M9_UM9_2_ParC7_PT3_line3, M9_UM9_2_ParC7_line3);
inv M9_UM9_2_ParC7_PT4_Xo3_0(M9_UM9_2_ParC7_line1, M9_UM9_2_ParC7_PT4_NotA);
inv M9_UM9_2_ParC7_PT4_Xo3_1(M9_UM9_2_ParC7_line2, M9_UM9_2_ParC7_PT4_NotB);
inv M9_UM9_2_ParC7_PT4_Xo3_2(M9_UM9_2_ParC7_line3, M9_UM9_2_ParC7_PT4_NotC);
and3 M9_UM9_2_ParC7_PT4_Xo3_3(M9_UM9_2_ParC7_PT4_NotA, M9_UM9_2_ParC7_PT4_NotB, M9_UM9_2_ParC7_line3, M9_UM9_2_ParC7_PT4_line3);
and3 M9_UM9_2_ParC7_PT4_Xo3_4(M9_UM9_2_ParC7_PT4_NotA, M9_UM9_2_ParC7_line2, M9_UM9_2_ParC7_PT4_NotC, M9_UM9_2_ParC7_PT4_line4);
and3 M9_UM9_2_ParC7_PT4_Xo3_5(M9_UM9_2_ParC7_line1, M9_UM9_2_ParC7_PT4_NotB, M9_UM9_2_ParC7_PT4_NotC, M9_UM9_2_ParC7_PT4_line5);
and3 M9_UM9_2_ParC7_PT4_Xo3_6(M9_UM9_2_ParC7_line1, M9_UM9_2_ParC7_line2, M9_UM9_2_ParC7_line3, M9_UM9_2_ParC7_PT4_line6);
nor2 M9_UM9_2_ParC7_PT4_Xo3_7(M9_UM9_2_ParC7_PT4_line3, M9_UM9_2_ParC7_PT4_line4, M9_UM9_2_ParC7_PT4_line7);
nor2 M9_UM9_2_ParC7_PT4_Xo3_8(M9_UM9_2_ParC7_PT4_line5, M9_UM9_2_ParC7_PT4_line6, M9_UM9_2_ParC7_PT4_line8);
nand2 M9_UM9_2_ParC7_PT4_Xo3_9(M9_UM9_2_ParC7_PT4_line7, M9_UM9_2_ParC7_PT4_line8, M9_UM9_2_ParC7_line4);
inv M9_UM9_2_ParC7_PT5_Xo0(M9_UM9_2_ParC7_line0, M9_UM9_2_ParC7_PT5_NotA);
inv M9_UM9_2_ParC7_PT5_Xo1(M9_UM9_2_ParC7_line4, M9_UM9_2_ParC7_PT5_NotB);
nand2 M9_UM9_2_ParC7_PT5_Xo2(M9_UM9_2_ParC7_PT5_NotA, M9_UM9_2_ParC7_line4, M9_UM9_2_ParC7_PT5_line2);
nand2 M9_UM9_2_ParC7_PT5_Xo3(M9_UM9_2_ParC7_PT5_NotB, M9_UM9_2_ParC7_line0, M9_UM9_2_ParC7_PT5_line3);
nand2 M9_UM9_2_ParC7_PT5_Xo4(M9_UM9_2_ParC7_PT5_line2, M9_UM9_2_ParC7_PT5_line3, M9_UM9_2_YaP3);
inv M9_UM9_2_ParC8_PT0_Xo0(YBbus_5, M9_UM9_2_ParC8_PT0_NotA);
inv M9_UM9_2_ParC8_PT0_Xo1(YBbus_6, M9_UM9_2_ParC8_PT0_NotB);
nand2 M9_UM9_2_ParC8_PT0_Xo2(M9_UM9_2_ParC8_PT0_NotA, YBbus_6, M9_UM9_2_ParC8_PT0_line2);
nand2 M9_UM9_2_ParC8_PT0_Xo3(M9_UM9_2_ParC8_PT0_NotB, YBbus_5, M9_UM9_2_ParC8_PT0_line3);
nand2 M9_UM9_2_ParC8_PT0_Xo4(M9_UM9_2_ParC8_PT0_line2, M9_UM9_2_ParC8_PT0_line3, M9_UM9_2_ParC8_line0);
inv M9_UM9_2_ParC8_PT1_Xo0(YBbus_7, M9_UM9_2_ParC8_PT1_NotA);
inv M9_UM9_2_ParC8_PT1_Xo1(YBbus_8, M9_UM9_2_ParC8_PT1_NotB);
nand2 M9_UM9_2_ParC8_PT1_Xo2(M9_UM9_2_ParC8_PT1_NotA, YBbus_8, M9_UM9_2_ParC8_PT1_line2);
nand2 M9_UM9_2_ParC8_PT1_Xo3(M9_UM9_2_ParC8_PT1_NotB, YBbus_7, M9_UM9_2_ParC8_PT1_line3);
nand2 M9_UM9_2_ParC8_PT1_Xo4(M9_UM9_2_ParC8_PT1_line2, M9_UM9_2_ParC8_PT1_line3, M9_UM9_2_ParC8_line1);
inv M9_UM9_2_ParC8_PT2_Xo0(YBbus_1, M9_UM9_2_ParC8_PT2_NotA);
inv M9_UM9_2_ParC8_PT2_Xo1(YBbus_2, M9_UM9_2_ParC8_PT2_NotB);
nand2 M9_UM9_2_ParC8_PT2_Xo2(M9_UM9_2_ParC8_PT2_NotA, YBbus_2, M9_UM9_2_ParC8_PT2_line2);
nand2 M9_UM9_2_ParC8_PT2_Xo3(M9_UM9_2_ParC8_PT2_NotB, YBbus_1, M9_UM9_2_ParC8_PT2_line3);
nand2 M9_UM9_2_ParC8_PT2_Xo4(M9_UM9_2_ParC8_PT2_line2, M9_UM9_2_ParC8_PT2_line3, M9_UM9_2_ParC8_line2);
inv M9_UM9_2_ParC8_PT3_Xo0(M9_UM9_1_PCYBtempbus_0, M9_UM9_2_ParC8_PT3_NotA);
inv M9_UM9_2_ParC8_PT3_Xo1(M9_UM9_1_PCYBtempbus_1, M9_UM9_2_ParC8_PT3_NotB);
nand2 M9_UM9_2_ParC8_PT3_Xo2(M9_UM9_2_ParC8_PT3_NotA, M9_UM9_1_PCYBtempbus_1, M9_UM9_2_ParC8_PT3_line2);
nand2 M9_UM9_2_ParC8_PT3_Xo3(M9_UM9_2_ParC8_PT3_NotB, M9_UM9_1_PCYBtempbus_0, M9_UM9_2_ParC8_PT3_line3);
nand2 M9_UM9_2_ParC8_PT3_Xo4(M9_UM9_2_ParC8_PT3_line2, M9_UM9_2_ParC8_PT3_line3, M9_UM9_2_ParC8_line3);
inv M9_UM9_2_ParC8_PT4_Xo0(YBbus_3, M9_UM9_2_ParC8_PT4_NotA);
inv M9_UM9_2_ParC8_PT4_Xo1(YBbus_4, M9_UM9_2_ParC8_PT4_NotB);
nand2 M9_UM9_2_ParC8_PT4_Xo2(M9_UM9_2_ParC8_PT4_NotA, YBbus_4, M9_UM9_2_ParC8_PT4_line2);
nand2 M9_UM9_2_ParC8_PT4_Xo3(M9_UM9_2_ParC8_PT4_NotB, YBbus_3, M9_UM9_2_ParC8_PT4_line3);
nand2 M9_UM9_2_ParC8_PT4_Xo4(M9_UM9_2_ParC8_PT4_line2, M9_UM9_2_ParC8_PT4_line3, M9_UM9_2_ParC8_line4);
inv M9_UM9_2_ParC8_PT5_Xo0(M9_UM9_2_ParC8_line0, M9_UM9_2_ParC8_PT5_NotA);
inv M9_UM9_2_ParC8_PT5_Xo1(M9_UM9_2_ParC8_line1, M9_UM9_2_ParC8_PT5_NotB);
nand2 M9_UM9_2_ParC8_PT5_Xo2(M9_UM9_2_ParC8_PT5_NotA, M9_UM9_2_ParC8_line1, M9_UM9_2_ParC8_PT5_line2);
nand2 M9_UM9_2_ParC8_PT5_Xo3(M9_UM9_2_ParC8_PT5_NotB, M9_UM9_2_ParC8_line0, M9_UM9_2_ParC8_PT5_line3);
nand2 M9_UM9_2_ParC8_PT5_Xo4(M9_UM9_2_ParC8_PT5_line2, M9_UM9_2_ParC8_PT5_line3, M9_UM9_2_ParC8_line5);
inv M9_UM9_2_ParC8_PT6_Xo3_0(M9_UM9_2_ParC8_line2, M9_UM9_2_ParC8_PT6_NotA);
inv M9_UM9_2_ParC8_PT6_Xo3_1(M9_UM9_2_ParC8_line3, M9_UM9_2_ParC8_PT6_NotB);
inv M9_UM9_2_ParC8_PT6_Xo3_2(M9_UM9_2_ParC8_line4, M9_UM9_2_ParC8_PT6_NotC);
and3 M9_UM9_2_ParC8_PT6_Xo3_3(M9_UM9_2_ParC8_PT6_NotA, M9_UM9_2_ParC8_PT6_NotB, M9_UM9_2_ParC8_line4, M9_UM9_2_ParC8_PT6_line3);
and3 M9_UM9_2_ParC8_PT6_Xo3_4(M9_UM9_2_ParC8_PT6_NotA, M9_UM9_2_ParC8_line3, M9_UM9_2_ParC8_PT6_NotC, M9_UM9_2_ParC8_PT6_line4);
and3 M9_UM9_2_ParC8_PT6_Xo3_5(M9_UM9_2_ParC8_line2, M9_UM9_2_ParC8_PT6_NotB, M9_UM9_2_ParC8_PT6_NotC, M9_UM9_2_ParC8_PT6_line5);
and3 M9_UM9_2_ParC8_PT6_Xo3_6(M9_UM9_2_ParC8_line2, M9_UM9_2_ParC8_line3, M9_UM9_2_ParC8_line4, M9_UM9_2_ParC8_PT6_line6);
nor2 M9_UM9_2_ParC8_PT6_Xo3_7(M9_UM9_2_ParC8_PT6_line3, M9_UM9_2_ParC8_PT6_line4, M9_UM9_2_ParC8_PT6_line7);
nor2 M9_UM9_2_ParC8_PT6_Xo3_8(M9_UM9_2_ParC8_PT6_line5, M9_UM9_2_ParC8_PT6_line6, M9_UM9_2_ParC8_PT6_line8);
nand2 M9_UM9_2_ParC8_PT6_Xo3_9(M9_UM9_2_ParC8_PT6_line7, M9_UM9_2_ParC8_PT6_line8, M9_UM9_2_ParC8_line6);
inv M9_UM9_2_ParC8_PT7_Xo0(M9_UM9_2_ParC8_line5, M9_UM9_2_ParC8_PT7_NotA);
inv M9_UM9_2_ParC8_PT7_Xo1(M9_UM9_2_ParC8_line6, M9_UM9_2_ParC8_PT7_NotB);
nand2 M9_UM9_2_ParC8_PT7_Xo2(M9_UM9_2_ParC8_PT7_NotA, M9_UM9_2_ParC8_line6, M9_UM9_2_ParC8_PT7_line2);
nand2 M9_UM9_2_ParC8_PT7_Xo3(M9_UM9_2_ParC8_PT7_NotB, M9_UM9_2_ParC8_line5, M9_UM9_2_ParC8_PT7_line3);
nand2 M9_UM9_2_ParC8_PT7_Xo4(M9_UM9_2_ParC8_PT7_line2, M9_UM9_2_ParC8_PT7_line3, M9_UM9_2_YbP0);
inv M9_UM9_2_ParC9_PT0_Xo0(YBbus_14, M9_UM9_2_ParC9_PT0_NotA);
inv M9_UM9_2_ParC9_PT0_Xo1(YBbus_15, M9_UM9_2_ParC9_PT0_NotB);
nand2 M9_UM9_2_ParC9_PT0_Xo2(M9_UM9_2_ParC9_PT0_NotA, YBbus_15, M9_UM9_2_ParC9_PT0_line2);
nand2 M9_UM9_2_ParC9_PT0_Xo3(M9_UM9_2_ParC9_PT0_NotB, YBbus_14, M9_UM9_2_ParC9_PT0_line3);
nand2 M9_UM9_2_ParC9_PT0_Xo4(M9_UM9_2_ParC9_PT0_line2, M9_UM9_2_ParC9_PT0_line3, M9_UM9_2_ParC9_line0);
inv M9_UM9_2_ParC9_PT1_Xo0(YBbus_16, M9_UM9_2_ParC9_PT1_NotA);
inv M9_UM9_2_ParC9_PT1_Xo1(YBbus_17, M9_UM9_2_ParC9_PT1_NotB);
nand2 M9_UM9_2_ParC9_PT1_Xo2(M9_UM9_2_ParC9_PT1_NotA, YBbus_17, M9_UM9_2_ParC9_PT1_line2);
nand2 M9_UM9_2_ParC9_PT1_Xo3(M9_UM9_2_ParC9_PT1_NotB, YBbus_16, M9_UM9_2_ParC9_PT1_line3);
nand2 M9_UM9_2_ParC9_PT1_Xo4(M9_UM9_2_ParC9_PT1_line2, M9_UM9_2_ParC9_PT1_line3, M9_UM9_2_ParC9_line1);
inv M9_UM9_2_ParC9_PT2_Xo0(YBbus_10, M9_UM9_2_ParC9_PT2_NotA);
inv M9_UM9_2_ParC9_PT2_Xo1(YBbus_11, M9_UM9_2_ParC9_PT2_NotB);
nand2 M9_UM9_2_ParC9_PT2_Xo2(M9_UM9_2_ParC9_PT2_NotA, YBbus_11, M9_UM9_2_ParC9_PT2_line2);
nand2 M9_UM9_2_ParC9_PT2_Xo3(M9_UM9_2_ParC9_PT2_NotB, YBbus_10, M9_UM9_2_ParC9_PT2_line3);
nand2 M9_UM9_2_ParC9_PT2_Xo4(M9_UM9_2_ParC9_PT2_line2, M9_UM9_2_ParC9_PT2_line3, M9_UM9_2_ParC9_line2);
inv M9_UM9_2_ParC9_PT3_Xo0(M9_UM9_1_PCYBtempbus_2, M9_UM9_2_ParC9_PT3_NotA);
inv M9_UM9_2_ParC9_PT3_Xo1(YBbus_9, M9_UM9_2_ParC9_PT3_NotB);
nand2 M9_UM9_2_ParC9_PT3_Xo2(M9_UM9_2_ParC9_PT3_NotA, YBbus_9, M9_UM9_2_ParC9_PT3_line2);
nand2 M9_UM9_2_ParC9_PT3_Xo3(M9_UM9_2_ParC9_PT3_NotB, M9_UM9_1_PCYBtempbus_2, M9_UM9_2_ParC9_PT3_line3);
nand2 M9_UM9_2_ParC9_PT3_Xo4(M9_UM9_2_ParC9_PT3_line2, M9_UM9_2_ParC9_PT3_line3, M9_UM9_2_ParC9_line3);
inv M9_UM9_2_ParC9_PT4_Xo0(YBbus_12, M9_UM9_2_ParC9_PT4_NotA);
inv M9_UM9_2_ParC9_PT4_Xo1(YBbus_13, M9_UM9_2_ParC9_PT4_NotB);
nand2 M9_UM9_2_ParC9_PT4_Xo2(M9_UM9_2_ParC9_PT4_NotA, YBbus_13, M9_UM9_2_ParC9_PT4_line2);
nand2 M9_UM9_2_ParC9_PT4_Xo3(M9_UM9_2_ParC9_PT4_NotB, YBbus_12, M9_UM9_2_ParC9_PT4_line3);
nand2 M9_UM9_2_ParC9_PT4_Xo4(M9_UM9_2_ParC9_PT4_line2, M9_UM9_2_ParC9_PT4_line3, M9_UM9_2_ParC9_line4);
inv M9_UM9_2_ParC9_PT5_Xo0(M9_UM9_2_ParC9_line0, M9_UM9_2_ParC9_PT5_NotA);
inv M9_UM9_2_ParC9_PT5_Xo1(M9_UM9_2_ParC9_line1, M9_UM9_2_ParC9_PT5_NotB);
nand2 M9_UM9_2_ParC9_PT5_Xo2(M9_UM9_2_ParC9_PT5_NotA, M9_UM9_2_ParC9_line1, M9_UM9_2_ParC9_PT5_line2);
nand2 M9_UM9_2_ParC9_PT5_Xo3(M9_UM9_2_ParC9_PT5_NotB, M9_UM9_2_ParC9_line0, M9_UM9_2_ParC9_PT5_line3);
nand2 M9_UM9_2_ParC9_PT5_Xo4(M9_UM9_2_ParC9_PT5_line2, M9_UM9_2_ParC9_PT5_line3, M9_UM9_2_ParC9_line5);
inv M9_UM9_2_ParC9_PT6_Xo3_0(M9_UM9_2_ParC9_line2, M9_UM9_2_ParC9_PT6_NotA);
inv M9_UM9_2_ParC9_PT6_Xo3_1(M9_UM9_2_ParC9_line3, M9_UM9_2_ParC9_PT6_NotB);
inv M9_UM9_2_ParC9_PT6_Xo3_2(M9_UM9_2_ParC9_line4, M9_UM9_2_ParC9_PT6_NotC);
and3 M9_UM9_2_ParC9_PT6_Xo3_3(M9_UM9_2_ParC9_PT6_NotA, M9_UM9_2_ParC9_PT6_NotB, M9_UM9_2_ParC9_line4, M9_UM9_2_ParC9_PT6_line3);
and3 M9_UM9_2_ParC9_PT6_Xo3_4(M9_UM9_2_ParC9_PT6_NotA, M9_UM9_2_ParC9_line3, M9_UM9_2_ParC9_PT6_NotC, M9_UM9_2_ParC9_PT6_line4);
and3 M9_UM9_2_ParC9_PT6_Xo3_5(M9_UM9_2_ParC9_line2, M9_UM9_2_ParC9_PT6_NotB, M9_UM9_2_ParC9_PT6_NotC, M9_UM9_2_ParC9_PT6_line5);
and3 M9_UM9_2_ParC9_PT6_Xo3_6(M9_UM9_2_ParC9_line2, M9_UM9_2_ParC9_line3, M9_UM9_2_ParC9_line4, M9_UM9_2_ParC9_PT6_line6);
nor2 M9_UM9_2_ParC9_PT6_Xo3_7(M9_UM9_2_ParC9_PT6_line3, M9_UM9_2_ParC9_PT6_line4, M9_UM9_2_ParC9_PT6_line7);
nor2 M9_UM9_2_ParC9_PT6_Xo3_8(M9_UM9_2_ParC9_PT6_line5, M9_UM9_2_ParC9_PT6_line6, M9_UM9_2_ParC9_PT6_line8);
nand2 M9_UM9_2_ParC9_PT6_Xo3_9(M9_UM9_2_ParC9_PT6_line7, M9_UM9_2_ParC9_PT6_line8, M9_UM9_2_ParC9_line6);
inv M9_UM9_2_ParC9_PT7_Xo0(M9_UM9_2_ParC9_line5, M9_UM9_2_ParC9_PT7_NotA);
inv M9_UM9_2_ParC9_PT7_Xo1(M9_UM9_2_ParC9_line6, M9_UM9_2_ParC9_PT7_NotB);
nand2 M9_UM9_2_ParC9_PT7_Xo2(M9_UM9_2_ParC9_PT7_NotA, M9_UM9_2_ParC9_line6, M9_UM9_2_ParC9_PT7_line2);
nand2 M9_UM9_2_ParC9_PT7_Xo3(M9_UM9_2_ParC9_PT7_NotB, M9_UM9_2_ParC9_line5, M9_UM9_2_ParC9_PT7_line3);
nand2 M9_UM9_2_ParC9_PT7_Xo4(M9_UM9_2_ParC9_PT7_line2, M9_UM9_2_ParC9_PT7_line3, M9_UM9_2_YbP1);
inv M9_UM9_2_ParC10_PT0_Xo0(YBbus_23, M9_UM9_2_ParC10_PT0_NotA);
inv M9_UM9_2_ParC10_PT0_Xo1(YBbus_24, M9_UM9_2_ParC10_PT0_NotB);
nand2 M9_UM9_2_ParC10_PT0_Xo2(M9_UM9_2_ParC10_PT0_NotA, YBbus_24, M9_UM9_2_ParC10_PT0_line2);
nand2 M9_UM9_2_ParC10_PT0_Xo3(M9_UM9_2_ParC10_PT0_NotB, YBbus_23, M9_UM9_2_ParC10_PT0_line3);
nand2 M9_UM9_2_ParC10_PT0_Xo4(M9_UM9_2_ParC10_PT0_line2, M9_UM9_2_ParC10_PT0_line3, M9_UM9_2_ParC10_line0);
inv M9_UM9_2_ParC10_PT1_Xo0(YBbus_25, M9_UM9_2_ParC10_PT1_NotA);
inv M9_UM9_2_ParC10_PT1_Xo1(YBbus_26, M9_UM9_2_ParC10_PT1_NotB);
nand2 M9_UM9_2_ParC10_PT1_Xo2(M9_UM9_2_ParC10_PT1_NotA, YBbus_26, M9_UM9_2_ParC10_PT1_line2);
nand2 M9_UM9_2_ParC10_PT1_Xo3(M9_UM9_2_ParC10_PT1_NotB, YBbus_25, M9_UM9_2_ParC10_PT1_line3);
nand2 M9_UM9_2_ParC10_PT1_Xo4(M9_UM9_2_ParC10_PT1_line2, M9_UM9_2_ParC10_PT1_line3, M9_UM9_2_ParC10_line1);
inv M9_UM9_2_ParC10_PT2_Xo0(YBbus_19, M9_UM9_2_ParC10_PT2_NotA);
inv M9_UM9_2_ParC10_PT2_Xo1(YBbus_20, M9_UM9_2_ParC10_PT2_NotB);
nand2 M9_UM9_2_ParC10_PT2_Xo2(M9_UM9_2_ParC10_PT2_NotA, YBbus_20, M9_UM9_2_ParC10_PT2_line2);
nand2 M9_UM9_2_ParC10_PT2_Xo3(M9_UM9_2_ParC10_PT2_NotB, YBbus_19, M9_UM9_2_ParC10_PT2_line3);
nand2 M9_UM9_2_ParC10_PT2_Xo4(M9_UM9_2_ParC10_PT2_line2, M9_UM9_2_ParC10_PT2_line3, M9_UM9_2_ParC10_line2);
inv M9_UM9_2_ParC10_PT3_Xo0(M9_UM9_1_PCYBtempbus_3, M9_UM9_2_ParC10_PT3_NotA);
inv M9_UM9_2_ParC10_PT3_Xo1(YBbus_18, M9_UM9_2_ParC10_PT3_NotB);
nand2 M9_UM9_2_ParC10_PT3_Xo2(M9_UM9_2_ParC10_PT3_NotA, YBbus_18, M9_UM9_2_ParC10_PT3_line2);
nand2 M9_UM9_2_ParC10_PT3_Xo3(M9_UM9_2_ParC10_PT3_NotB, M9_UM9_1_PCYBtempbus_3, M9_UM9_2_ParC10_PT3_line3);
nand2 M9_UM9_2_ParC10_PT3_Xo4(M9_UM9_2_ParC10_PT3_line2, M9_UM9_2_ParC10_PT3_line3, M9_UM9_2_ParC10_line3);
inv M9_UM9_2_ParC10_PT4_Xo0(YBbus_21, M9_UM9_2_ParC10_PT4_NotA);
inv M9_UM9_2_ParC10_PT4_Xo1(YBbus_22, M9_UM9_2_ParC10_PT4_NotB);
nand2 M9_UM9_2_ParC10_PT4_Xo2(M9_UM9_2_ParC10_PT4_NotA, YBbus_22, M9_UM9_2_ParC10_PT4_line2);
nand2 M9_UM9_2_ParC10_PT4_Xo3(M9_UM9_2_ParC10_PT4_NotB, YBbus_21, M9_UM9_2_ParC10_PT4_line3);
nand2 M9_UM9_2_ParC10_PT4_Xo4(M9_UM9_2_ParC10_PT4_line2, M9_UM9_2_ParC10_PT4_line3, M9_UM9_2_ParC10_line4);
inv M9_UM9_2_ParC10_PT5_Xo0(M9_UM9_2_ParC10_line0, M9_UM9_2_ParC10_PT5_NotA);
inv M9_UM9_2_ParC10_PT5_Xo1(M9_UM9_2_ParC10_line1, M9_UM9_2_ParC10_PT5_NotB);
nand2 M9_UM9_2_ParC10_PT5_Xo2(M9_UM9_2_ParC10_PT5_NotA, M9_UM9_2_ParC10_line1, M9_UM9_2_ParC10_PT5_line2);
nand2 M9_UM9_2_ParC10_PT5_Xo3(M9_UM9_2_ParC10_PT5_NotB, M9_UM9_2_ParC10_line0, M9_UM9_2_ParC10_PT5_line3);
nand2 M9_UM9_2_ParC10_PT5_Xo4(M9_UM9_2_ParC10_PT5_line2, M9_UM9_2_ParC10_PT5_line3, M9_UM9_2_ParC10_line5);
inv M9_UM9_2_ParC10_PT6_Xo3_0(M9_UM9_2_ParC10_line2, M9_UM9_2_ParC10_PT6_NotA);
inv M9_UM9_2_ParC10_PT6_Xo3_1(M9_UM9_2_ParC10_line3, M9_UM9_2_ParC10_PT6_NotB);
inv M9_UM9_2_ParC10_PT6_Xo3_2(M9_UM9_2_ParC10_line4, M9_UM9_2_ParC10_PT6_NotC);
and3 M9_UM9_2_ParC10_PT6_Xo3_3(M9_UM9_2_ParC10_PT6_NotA, M9_UM9_2_ParC10_PT6_NotB, M9_UM9_2_ParC10_line4, M9_UM9_2_ParC10_PT6_line3);
and3 M9_UM9_2_ParC10_PT6_Xo3_4(M9_UM9_2_ParC10_PT6_NotA, M9_UM9_2_ParC10_line3, M9_UM9_2_ParC10_PT6_NotC, M9_UM9_2_ParC10_PT6_line4);
and3 M9_UM9_2_ParC10_PT6_Xo3_5(M9_UM9_2_ParC10_line2, M9_UM9_2_ParC10_PT6_NotB, M9_UM9_2_ParC10_PT6_NotC, M9_UM9_2_ParC10_PT6_line5);
and3 M9_UM9_2_ParC10_PT6_Xo3_6(M9_UM9_2_ParC10_line2, M9_UM9_2_ParC10_line3, M9_UM9_2_ParC10_line4, M9_UM9_2_ParC10_PT6_line6);
nor2 M9_UM9_2_ParC10_PT6_Xo3_7(M9_UM9_2_ParC10_PT6_line3, M9_UM9_2_ParC10_PT6_line4, M9_UM9_2_ParC10_PT6_line7);
nor2 M9_UM9_2_ParC10_PT6_Xo3_8(M9_UM9_2_ParC10_PT6_line5, M9_UM9_2_ParC10_PT6_line6, M9_UM9_2_ParC10_PT6_line8);
nand2 M9_UM9_2_ParC10_PT6_Xo3_9(M9_UM9_2_ParC10_PT6_line7, M9_UM9_2_ParC10_PT6_line8, M9_UM9_2_ParC10_line6);
inv M9_UM9_2_ParC10_PT7_Xo0(M9_UM9_2_ParC10_line5, M9_UM9_2_ParC10_PT7_NotA);
inv M9_UM9_2_ParC10_PT7_Xo1(M9_UM9_2_ParC10_line6, M9_UM9_2_ParC10_PT7_NotB);
nand2 M9_UM9_2_ParC10_PT7_Xo2(M9_UM9_2_ParC10_PT7_NotA, M9_UM9_2_ParC10_line6, M9_UM9_2_ParC10_PT7_line2);
nand2 M9_UM9_2_ParC10_PT7_Xo3(M9_UM9_2_ParC10_PT7_NotB, M9_UM9_2_ParC10_line5, M9_UM9_2_ParC10_PT7_line3);
nand2 M9_UM9_2_ParC10_PT7_Xo4(M9_UM9_2_ParC10_PT7_line2, M9_UM9_2_ParC10_PT7_line3, M9_UM9_2_YbP2);
inv M9_UM9_2_ParC11_PT0_Xo0(M9_PCYBbus_4, M9_UM9_2_ParC11_PT0_NotA);
inv M9_UM9_2_ParC11_PT0_Xo1(M9_PCYBbus_5, M9_UM9_2_ParC11_PT0_NotB);
nand2 M9_UM9_2_ParC11_PT0_Xo2(M9_UM9_2_ParC11_PT0_NotA, M9_PCYBbus_5, M9_UM9_2_ParC11_PT0_line2);
nand2 M9_UM9_2_ParC11_PT0_Xo3(M9_UM9_2_ParC11_PT0_NotB, M9_PCYBbus_4, M9_UM9_2_ParC11_PT0_line3);
nand2 M9_UM9_2_ParC11_PT0_Xo4(M9_UM9_2_ParC11_PT0_line2, M9_UM9_2_ParC11_PT0_line3, M9_UM9_2_ParC11_line0);
inv M9_UM9_2_ParC11_PT1_Xo0(M9_PCYBbus_6, M9_UM9_2_ParC11_PT1_NotA);
inv M9_UM9_2_ParC11_PT1_Xo1(YBbus_27, M9_UM9_2_ParC11_PT1_NotB);
nand2 M9_UM9_2_ParC11_PT1_Xo2(M9_UM9_2_ParC11_PT1_NotA, YBbus_27, M9_UM9_2_ParC11_PT1_line2);
nand2 M9_UM9_2_ParC11_PT1_Xo3(M9_UM9_2_ParC11_PT1_NotB, M9_PCYBbus_6, M9_UM9_2_ParC11_PT1_line3);
nand2 M9_UM9_2_ParC11_PT1_Xo4(M9_UM9_2_ParC11_PT1_line2, M9_UM9_2_ParC11_PT1_line3, M9_UM9_2_ParC11_line1);
inv M9_UM9_2_ParC11_PT2_Xo0(YBbus_28, M9_UM9_2_ParC11_PT2_NotA);
inv M9_UM9_2_ParC11_PT2_Xo1(YBbus_29, M9_UM9_2_ParC11_PT2_NotB);
nand2 M9_UM9_2_ParC11_PT2_Xo2(M9_UM9_2_ParC11_PT2_NotA, YBbus_29, M9_UM9_2_ParC11_PT2_line2);
nand2 M9_UM9_2_ParC11_PT2_Xo3(M9_UM9_2_ParC11_PT2_NotB, YBbus_28, M9_UM9_2_ParC11_PT2_line3);
nand2 M9_UM9_2_ParC11_PT2_Xo4(M9_UM9_2_ParC11_PT2_line2, M9_UM9_2_ParC11_PT2_line3, M9_UM9_2_ParC11_line2);
inv M9_UM9_2_ParC11_PT3_Xo0(YBbus_30, M9_UM9_2_ParC11_PT3_NotA);
inv M9_UM9_2_ParC11_PT3_Xo1(YBbus_31, M9_UM9_2_ParC11_PT3_NotB);
nand2 M9_UM9_2_ParC11_PT3_Xo2(M9_UM9_2_ParC11_PT3_NotA, YBbus_31, M9_UM9_2_ParC11_PT3_line2);
nand2 M9_UM9_2_ParC11_PT3_Xo3(M9_UM9_2_ParC11_PT3_NotB, YBbus_30, M9_UM9_2_ParC11_PT3_line3);
nand2 M9_UM9_2_ParC11_PT3_Xo4(M9_UM9_2_ParC11_PT3_line2, M9_UM9_2_ParC11_PT3_line3, M9_UM9_2_ParC11_line3);
inv M9_UM9_2_ParC11_PT4_Xo3_0(M9_UM9_2_ParC11_line1, M9_UM9_2_ParC11_PT4_NotA);
inv M9_UM9_2_ParC11_PT4_Xo3_1(M9_UM9_2_ParC11_line2, M9_UM9_2_ParC11_PT4_NotB);
inv M9_UM9_2_ParC11_PT4_Xo3_2(M9_UM9_2_ParC11_line3, M9_UM9_2_ParC11_PT4_NotC);
and3 M9_UM9_2_ParC11_PT4_Xo3_3(M9_UM9_2_ParC11_PT4_NotA, M9_UM9_2_ParC11_PT4_NotB, M9_UM9_2_ParC11_line3, M9_UM9_2_ParC11_PT4_line3);
and3 M9_UM9_2_ParC11_PT4_Xo3_4(M9_UM9_2_ParC11_PT4_NotA, M9_UM9_2_ParC11_line2, M9_UM9_2_ParC11_PT4_NotC, M9_UM9_2_ParC11_PT4_line4);
and3 M9_UM9_2_ParC11_PT4_Xo3_5(M9_UM9_2_ParC11_line1, M9_UM9_2_ParC11_PT4_NotB, M9_UM9_2_ParC11_PT4_NotC, M9_UM9_2_ParC11_PT4_line5);
and3 M9_UM9_2_ParC11_PT4_Xo3_6(M9_UM9_2_ParC11_line1, M9_UM9_2_ParC11_line2, M9_UM9_2_ParC11_line3, M9_UM9_2_ParC11_PT4_line6);
nor2 M9_UM9_2_ParC11_PT4_Xo3_7(M9_UM9_2_ParC11_PT4_line3, M9_UM9_2_ParC11_PT4_line4, M9_UM9_2_ParC11_PT4_line7);
nor2 M9_UM9_2_ParC11_PT4_Xo3_8(M9_UM9_2_ParC11_PT4_line5, M9_UM9_2_ParC11_PT4_line6, M9_UM9_2_ParC11_PT4_line8);
nand2 M9_UM9_2_ParC11_PT4_Xo3_9(M9_UM9_2_ParC11_PT4_line7, M9_UM9_2_ParC11_PT4_line8, M9_UM9_2_ParC11_line4);
inv M9_UM9_2_ParC11_PT5_Xo0(M9_UM9_2_ParC11_line0, M9_UM9_2_ParC11_PT5_NotA);
inv M9_UM9_2_ParC11_PT5_Xo1(M9_UM9_2_ParC11_line4, M9_UM9_2_ParC11_PT5_NotB);
nand2 M9_UM9_2_ParC11_PT5_Xo2(M9_UM9_2_ParC11_PT5_NotA, M9_UM9_2_ParC11_line4, M9_UM9_2_ParC11_PT5_line2);
nand2 M9_UM9_2_ParC11_PT5_Xo3(M9_UM9_2_ParC11_PT5_NotB, M9_UM9_2_ParC11_line0, M9_UM9_2_ParC11_PT5_line3);
nand2 M9_UM9_2_ParC11_PT5_Xo4(M9_UM9_2_ParC11_PT5_line2, M9_UM9_2_ParC11_PT5_line3, M9_UM9_2_YbP3);
and4 M9_UM9_2_ParC12(M9_UM9_2_XaP0, M9_UM9_2_XaP1, M9_UM9_2_XaP2, M9_UM9_2_XaP3, M9_UM9_2_XaP);
and4 M9_UM9_2_ParC13(M9_UM9_2_YaP0, M9_UM9_2_YaP1, M9_UM9_2_YaP2, M9_UM9_2_YaP3, M9_UM9_2_YaP);
and4 M9_UM9_2_ParC14(M9_UM9_2_YbP0, M9_UM9_2_YbP1, M9_UM9_2_YbP2, M9_UM9_2_YbP3, M9_UM9_2_YbP);
and3 M9_UM9_2_ParC15(M9_UM9_2_XaP, M9_UM9_2_YaP, M9_UM9_2_YbP, M9_UM9_2_XYabP);
and3 M9_UM9_2_ParC16(M9_StrobeK0_1, M9_StrobeK2_3, M9_UM9_2_XYabP, M9_UM9_2_NotPar0);
inv M9_UM9_2_ParC17(M9_UM9_2_NotPar0, out418);
inv M9_UM9_2_ParC18(M9_UM9_2_XaP, out412);
inv M9_UM9_2_ParC19(M9_UM9_2_YaP, out414);
inv M9_UM9_2_ParC20(M9_UM9_2_YbP, out416);
buffer M10_Buf34_0_Buf8_0_Buf4_0(in3701, out542);
buffer M10_Buf34_0_Buf8_0_Buf4_1(in3705, out558);
buffer M10_Buf34_0_Buf8_0_Buf4_2(in3711, out556);
buffer M10_Buf34_0_Buf8_0_Buf4_3(in3717, out554);
buffer M10_Buf34_0_Buf8_1_Buf4_0(in3723, out552);
buffer M10_Buf34_0_Buf8_1_Buf4_1(in3729, out550);
buffer M10_Buf34_0_Buf8_1_Buf4_2(in3737, out548);
buffer M10_Buf34_0_Buf8_1_Buf4_3(in3743, out546);
buffer M10_Buf34_1_Buf8_0_Buf4_0(in3749, out544);
buffer M10_Buf34_1_Buf8_0_Buf4_1(in4394, out522);
buffer M10_Buf34_1_Buf8_0_Buf4_2(in4400, out538);
buffer M10_Buf34_1_Buf8_0_Buf4_3(in4405, out536);
buffer M10_Buf34_1_Buf8_1_Buf4_0(in4410, out534);
buffer M10_Buf34_1_Buf8_1_Buf4_1(in4415, out532);
buffer M10_Buf34_1_Buf8_1_Buf4_2(in4420, out530);
buffer M10_Buf34_1_Buf8_1_Buf4_3(in4427, out528);
buffer M10_Buf34_2_Buf8_0_Buf4_0(in4432, out526);
buffer M10_Buf34_2_Buf8_0_Buf4_1(in4437, out524);
buffer M10_Buf34_2_Buf8_0_Buf4_2(in2211, out478);
buffer M10_Buf34_2_Buf8_0_Buf4_3(in2218, out494);
buffer M10_Buf34_2_Buf8_1_Buf4_0(in2224, out492);
buffer M10_Buf34_2_Buf8_1_Buf4_1(in2230, out490);
buffer M10_Buf34_2_Buf8_1_Buf4_2(in2236, out488);
buffer M10_Buf34_2_Buf8_1_Buf4_3(in2239, out486);
buffer M10_Buf34_3_Buf8_0_Buf4_0(in2247, out484);
buffer M10_Buf34_3_Buf8_0_Buf4_1(in2253, out482);
buffer M10_Buf34_3_Buf8_0_Buf4_2(in2256, out480);
buffer M10_Buf34_3_Buf8_0_Buf4_3(in1462, out436);
buffer M10_Buf34_3_Buf8_1_Buf4_0(in1469, out448);
buffer M10_Buf34_3_Buf8_1_Buf4_1(in106, out446);
buffer M10_Buf34_3_Buf8_1_Buf4_2(in1480, out444);
buffer M10_Buf34_3_Buf8_1_Buf4_3(in1486, out442);
buffer M10_Buf34_4(in1492, out440);
buffer M10_Buf34_5(in1496, out438);
buffer M11_Buf4_0(in3698, out560);
buffer M11_Buf4_1(in4393, out540);
buffer M11_Buf4_2(in2208, out496);
buffer M11_Buf4_3(in1459, out450);
buffer M12_UM12_0(in1, out2);
and2 M12_UM12_1(in1, in163, out278);
inv M12_UM12_2(in15, out279);
and2 M12_UM12_3(in134, in133, M12_line3);
inv M12_UM12_4(in5, M12_line4);
nand2 M12_UM12_5(M12_line3, M12_line4, out292);
nand2 M12_UM12_6(in1197, M12_line4, out289);
inv M12_UM12_7(in57, M12_line7);
nand2 M12_UM12_8(M12_line7, M12_line4, out402);

assign out419 = out471;
assign out422 = out469;
assign out270 = CarryXbus_33;
assign out246 = CarryXbus_33;
assign out276 = out273;
assign out258 = M8_CarryOutYbus_33;
assign out264 = M8_CarryOutYbus_33;
assign out3 = out2;
assign out432 = out2;
assign out453 = out2;
assign out286 = out279;
assign out341 = out279;
assign out281 = out292;
assign out284 = out289;
assign out339 = in339;
assign vdd = 1'b1;
assign gnd = 1'b0;

endmodule
