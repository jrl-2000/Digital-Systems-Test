
//Verilog file of module c2670


`timescale 1 ns / 1ns

module c2670_net(G1,
G10,
G100,
G101,
G102,
G103,
G104,
G105,
G106,
G107,
G108,
G109,
G11,
G110,
G111,
G112,
G113,
G114,
G115,
G116,
G117,
G118,
G119,
G12,
G120,
G121,
G122,
G123,
G124,
G125,
G126,
G127,
G128,
G129,
G13,
G130,
G131,
G132,
G133,
G134,
G135,
G136,
G137,
G138,
G139,
G14,
G140,
G141,
G142,
G143,
G144,
G145,
G146,
G147,
G148,
G149,
G15,
G150,
G151,
G152,
G153,
G154,
G155,
G156,
G157,
G16,
G17,
G18,
G19,
G2,
G20,
G21,
G22,
G23,
G24,
G25,
G2531,
G2532,
G2533,
G2534,
G2535,
G2536,
G2537,
G2538,
G2539,
G2540,
G2541,
G2542,
G2543,
G2544,
G2545,
G2546,
G2547,
G2548,
G2549,
G2550,
G2551,
G2552,
G2553,
G2554,
G2555,
G2556,
G2557,
G2558,
G2559,
G2560,
G2561,
G2562,
G2563,
G2564,
G2565,
G2566,
G2567,
G2568,
G2569,
G2570,
G2571,
G2572,
G2573,
G2574,
G2575,
G2576,
G2577,
G2578,
G2579,
G2580,
G2581,
G2582,
G2583,
G2584,
G2585,
G2586,
G2587,
G2588,
G2589,
G2590,
G2591,
G2592,
G2593,
G2594,
G26,
G27,
G28,
G29,
G3,
G30,
G31,
G32,
G33,
G34,
G35,
G36,
G37,
G38,
G39,
G4,
G40,
G41,
G42,
G43,
G44,
G45,
G46,
G47,
G48,
G49,
G5,
G50,
G51,
G52,
G53,
G54,
G55,
G56,
G57,
G58,
G59,
G6,
G60,
G61,
G62,
G63,
G64,
G65,
G66,
G67,
G68,
G69,
G7,
G70,
G71,
G72,
G73,
G74,
G75,
G76,
G77,
G78,
G79,
G8,
G80,
G81,
G82,
G83,
G84,
G85,
G86,
G87,
G88,
G89,
G9,
G90,
G91,
G92,
G93,
G94,
G95,
G96,
G97,
G98,
G99);
input G1;
input G2;
input G3;
input G4;
input G5;
input G6;
input G7;
input G8;
input G9;
input G10;
input G11;
input G12;
input G13;
input G14;
input G15;
input G16;
input G17;
input G18;
input G19;
input G20;
input G21;
input G22;
input G23;
input G24;
input G25;
input G26;
input G27;
input G28;
input G29;
input G30;
input G31;
input G32;
input G33;
input G34;
input G35;
input G36;
input G37;
input G38;
input G39;
input G40;
input G41;
input G42;
input G43;
input G44;
input G45;
input G46;
input G47;
input G48;
input G49;
input G50;
input G51;
input G52;
input G53;
input G54;
input G55;
input G56;
input G57;
input G58;
input G59;
input G60;
input G61;
input G62;
input G63;
input G64;
input G65;
input G66;
input G67;
input G68;
input G69;
input G70;
input G71;
input G72;
input G73;
input G74;
input G75;
input G76;
input G77;
input G78;
input G79;
input G80;
input G81;
input G82;
input G83;
input G84;
input G85;
input G86;
input G87;
input G88;
input G89;
input G90;
input G91;
input G92;
input G93;
input G94;
input G95;
input G96;
input G97;
input G98;
input G99;
input G100;
input G101;
input G102;
input G103;
input G104;
input G105;
input G106;
input G107;
input G108;
input G109;
input G110;
input G111;
input G112;
input G113;
input G114;
input G115;
input G116;
input G117;
input G118;
input G119;
input G120;
input G121;
input G122;
input G123;
input G124;
input G125;
input G126;
input G127;
input G128;
input G129;
input G130;
input G131;
input G132;
input G133;
input G134;
input G135;
input G136;
input G137;
input G138;
input G139;
input G140;
input G141;
input G142;
input G143;
input G144;
input G145;
input G146;
input G147;
input G148;
input G149;
input G150;
input G151;
input G152;
input G153;
input G154;
input G155;
input G156;
input G157;

output G2531;
output G2532;
output G2533;
output G2534;
output G2535;
output G2536;
output G2537;
output G2538;
output G2539;
output G2540;
output G2541;
output G2542;
output G2543;
output G2544;
output G2545;
output G2546;
output G2547;
output G2548;
output G2549;
output G2550;
output G2551;
output G2552;
output G2553;
output G2554;
output G2555;
output G2556;
output G2557;
output G2558;
output G2559;
output G2560;
output G2561;
output G2562;
output G2563;
output G2564;
output G2565;
output G2566;
output G2567;
output G2568;
output G2569;
output G2570;
output G2571;
output G2572;
output G2573;
output G2574;
output G2575;
output G2576;
output G2577;
output G2578;
output G2579;
output G2580;
output G2581;
output G2582;
output G2583;
output G2584;
output G2585;
output G2586;
output G2587;
output G2588;
output G2589;
output G2590;
output G2591;
output G2592;
output G2593;
output G2594;

wire
c2670_wire_1,
c2670_wire_2,
c2670_wire_3,
c2670_wire_4,
c2670_wire_5,
c2670_wire_6,
c2670_wire_7,
c2670_wire_8,
c2670_wire_9,
c2670_wire_10,
c2670_wire_11,
c2670_wire_12,
c2670_wire_13,
c2670_wire_14,
c2670_wire_15,
c2670_wire_16,
c2670_wire_17,
c2670_wire_18,
c2670_wire_19,
c2670_wire_20,
c2670_wire_21,
c2670_wire_22,
c2670_wire_23,
c2670_wire_24,
c2670_wire_25,
c2670_wire_26,
c2670_wire_27,
c2670_wire_28,
c2670_wire_29,
c2670_wire_30,
c2670_wire_31,
c2670_wire_32,
c2670_wire_33,
c2670_wire_34,
c2670_wire_35,
c2670_wire_36,
c2670_wire_37,
c2670_wire_38,
c2670_wire_39,
c2670_wire_40,
c2670_wire_41,
c2670_wire_42,
c2670_wire_43,
c2670_wire_44,
c2670_wire_45,
c2670_wire_46,
c2670_wire_47,
c2670_wire_48,
c2670_wire_49,
c2670_wire_50,
c2670_wire_51,
c2670_wire_52,
c2670_wire_53,
c2670_wire_54,
c2670_wire_55,
c2670_wire_56,
c2670_wire_57,
c2670_wire_58,
c2670_wire_59,
c2670_wire_60,
c2670_wire_61,
c2670_wire_62,
c2670_wire_63,
c2670_wire_64,
c2670_wire_65,
c2670_wire_66,
c2670_wire_67,
c2670_wire_68,
c2670_wire_69,
c2670_wire_70,
c2670_wire_71,
c2670_wire_72,
c2670_wire_73,
c2670_wire_74,
c2670_wire_75,
c2670_wire_76,
c2670_wire_77,
c2670_wire_78,
c2670_wire_79,
c2670_wire_80,
c2670_wire_81,
c2670_wire_82,
c2670_wire_83,
c2670_wire_84,
c2670_wire_85,
c2670_wire_86,
c2670_wire_87,
c2670_wire_88,
c2670_wire_89,
c2670_wire_90,
c2670_wire_91,
c2670_wire_92,
c2670_wire_93,
c2670_wire_94,
c2670_wire_95,
c2670_wire_96,
c2670_wire_97,
c2670_wire_98,
c2670_wire_99,
c2670_wire_100,
c2670_wire_101,
c2670_wire_102,
c2670_wire_103,
c2670_wire_104,
c2670_wire_105,
c2670_wire_106,
c2670_wire_107,
c2670_wire_108,
c2670_wire_109,
c2670_wire_110,
c2670_wire_111,
c2670_wire_112,
c2670_wire_113,
c2670_wire_114,
c2670_wire_115,
c2670_wire_116,
c2670_wire_117,
c2670_wire_118,
c2670_wire_119,
c2670_wire_120,
c2670_wire_121,
c2670_wire_122,
c2670_wire_123,
c2670_wire_124,
c2670_wire_125,
c2670_wire_126,
c2670_wire_127,
c2670_wire_128,
c2670_wire_129,
c2670_wire_130,
c2670_wire_131,
c2670_wire_132,
c2670_wire_133,
c2670_wire_134,
c2670_wire_135,
c2670_wire_136,
c2670_wire_137,
c2670_wire_138,
c2670_wire_139,
c2670_wire_140,
c2670_wire_141,
c2670_wire_142,
c2670_wire_143,
c2670_wire_144,
c2670_wire_145,
c2670_wire_146,
c2670_wire_147,
c2670_wire_148,
c2670_wire_149,
c2670_wire_150,
c2670_wire_151,
c2670_wire_152,
c2670_wire_153,
c2670_wire_154,
c2670_wire_155,
c2670_wire_156,
c2670_wire_157,
c2670_wire_158,
c2670_wire_159,
c2670_wire_160,
c2670_wire_161,
c2670_wire_162,
c2670_wire_163,
c2670_wire_164,
c2670_wire_165,
c2670_wire_166,
c2670_wire_167,
c2670_wire_168,
c2670_wire_169,
c2670_wire_170,
c2670_wire_171,
c2670_wire_172,
c2670_wire_173,
c2670_wire_174,
c2670_wire_175,
c2670_wire_176,
c2670_wire_177,
c2670_wire_178,
c2670_wire_179,
c2670_wire_180,
c2670_wire_181,
c2670_wire_182,
c2670_wire_183,
c2670_wire_184,
c2670_wire_185,
c2670_wire_186,
c2670_wire_187,
c2670_wire_188,
c2670_wire_189,
c2670_wire_190,
c2670_wire_191,
c2670_wire_192,
c2670_wire_193,
c2670_wire_194,
c2670_wire_195,
c2670_wire_196,
c2670_wire_197,
c2670_wire_198,
c2670_wire_199,
c2670_wire_200,
c2670_wire_201,
c2670_wire_202,
c2670_wire_203,
c2670_wire_204,
c2670_wire_205,
c2670_wire_206,
c2670_wire_207,
c2670_wire_208,
c2670_wire_209,
c2670_wire_210,
c2670_wire_211,
c2670_wire_212,
c2670_wire_213,
c2670_wire_214,
c2670_wire_215,
c2670_wire_216,
c2670_wire_217,
c2670_wire_218,
c2670_wire_219,
c2670_wire_220,
c2670_wire_221,
c2670_wire_222,
c2670_wire_223,
c2670_wire_224,
c2670_wire_225,
c2670_wire_226,
c2670_wire_227,
c2670_wire_228,
c2670_wire_229,
c2670_wire_230,
c2670_wire_231,
c2670_wire_232,
c2670_wire_233,
c2670_wire_234,
c2670_wire_235,
c2670_wire_236,
c2670_wire_237,
c2670_wire_238,
c2670_wire_239,
c2670_wire_240,
c2670_wire_241,
c2670_wire_242,
c2670_wire_243,
c2670_wire_244,
c2670_wire_245,
c2670_wire_246,
c2670_wire_247,
c2670_wire_248,
c2670_wire_249,
c2670_wire_250,
c2670_wire_251,
c2670_wire_252,
c2670_wire_253,
c2670_wire_254,
c2670_wire_255,
c2670_wire_256,
c2670_wire_257,
c2670_wire_258,
c2670_wire_259,
c2670_wire_260,
c2670_wire_261,
c2670_wire_262,
c2670_wire_263,
c2670_wire_264,
c2670_wire_265,
c2670_wire_266,
c2670_wire_267,
c2670_wire_268,
c2670_wire_269,
c2670_wire_270,
c2670_wire_271,
c2670_wire_272,
c2670_wire_273,
c2670_wire_274,
c2670_wire_275,
c2670_wire_276,
c2670_wire_277,
c2670_wire_278,
c2670_wire_279,
c2670_wire_280,
c2670_wire_281,
c2670_wire_282,
c2670_wire_283,
c2670_wire_284,
c2670_wire_285,
c2670_wire_286,
c2670_wire_287,
c2670_wire_288,
c2670_wire_289,
c2670_wire_290,
c2670_wire_291,
c2670_wire_292,
c2670_wire_293,
c2670_wire_294,
c2670_wire_295,
c2670_wire_296,
c2670_wire_297,
c2670_wire_298,
c2670_wire_299,
c2670_wire_300,
c2670_wire_301,
c2670_wire_302,
c2670_wire_303,
c2670_wire_304,
c2670_wire_305,
c2670_wire_306,
c2670_wire_307,
c2670_wire_308,
c2670_wire_309,
c2670_wire_310,
c2670_wire_311,
c2670_wire_312,
c2670_wire_313,
c2670_wire_314,
c2670_wire_315,
c2670_wire_316,
c2670_wire_317,
c2670_wire_318,
c2670_wire_319,
c2670_wire_320,
c2670_wire_321,
c2670_wire_322,
c2670_wire_323,
c2670_wire_324,
c2670_wire_325,
c2670_wire_326,
c2670_wire_327,
c2670_wire_328,
c2670_wire_329,
c2670_wire_330,
c2670_wire_331,
c2670_wire_332,
c2670_wire_333,
c2670_wire_334,
c2670_wire_335,
c2670_wire_336,
c2670_wire_337,
c2670_wire_338,
c2670_wire_339,
c2670_wire_340,
c2670_wire_341,
c2670_wire_342,
c2670_wire_343,
c2670_wire_344,
c2670_wire_345,
c2670_wire_346,
c2670_wire_347,
c2670_wire_348,
c2670_wire_349,
c2670_wire_350,
c2670_wire_351,
c2670_wire_352,
c2670_wire_353,
c2670_wire_354,
c2670_wire_355,
c2670_wire_356,
c2670_wire_357,
c2670_wire_358,
c2670_wire_359,
c2670_wire_360,
c2670_wire_361,
c2670_wire_362,
c2670_wire_363,
c2670_wire_364,
c2670_wire_365,
c2670_wire_366,
c2670_wire_367,
c2670_wire_368,
c2670_wire_369,
c2670_wire_370,
c2670_wire_371,
c2670_wire_372,
c2670_wire_373,
c2670_wire_374,
c2670_wire_375,
c2670_wire_376,
c2670_wire_377,
c2670_wire_378,
c2670_wire_379,
c2670_wire_380,
c2670_wire_381,
c2670_wire_382,
c2670_wire_383,
c2670_wire_384,
c2670_wire_385,
c2670_wire_386,
c2670_wire_387,
c2670_wire_388,
c2670_wire_389,
c2670_wire_390,
c2670_wire_391,
c2670_wire_392,
c2670_wire_393,
c2670_wire_394,
c2670_wire_395,
c2670_wire_396,
c2670_wire_397,
c2670_wire_398,
c2670_wire_399,
c2670_wire_400,
c2670_wire_401,
c2670_wire_402,
c2670_wire_403,
c2670_wire_404,
c2670_wire_405,
c2670_wire_406,
c2670_wire_407,
c2670_wire_408,
c2670_wire_409,
c2670_wire_410,
c2670_wire_411,
c2670_wire_412,
c2670_wire_413,
c2670_wire_414,
c2670_wire_415,
c2670_wire_416,
c2670_wire_417,
c2670_wire_418,
c2670_wire_419,
c2670_wire_420,
c2670_wire_421,
c2670_wire_422,
c2670_wire_423,
c2670_wire_424,
c2670_wire_425,
c2670_wire_426,
c2670_wire_427,
c2670_wire_428,
c2670_wire_429,
c2670_wire_430,
c2670_wire_431,
c2670_wire_432,
c2670_wire_433,
c2670_wire_434,
c2670_wire_435,
c2670_wire_436,
c2670_wire_437,
c2670_wire_438,
c2670_wire_439,
c2670_wire_440,
c2670_wire_441,
c2670_wire_442,
c2670_wire_443,
c2670_wire_444,
c2670_wire_445,
c2670_wire_446,
c2670_wire_447,
c2670_wire_448,
c2670_wire_449,
c2670_wire_450,
c2670_wire_451,
c2670_wire_452,
c2670_wire_453,
c2670_wire_454,
c2670_wire_455,
c2670_wire_456,
c2670_wire_457,
c2670_wire_458,
c2670_wire_459,
c2670_wire_460,
c2670_wire_461,
c2670_wire_462,
c2670_wire_463,
c2670_wire_464,
c2670_wire_465,
c2670_wire_466,
c2670_wire_467,
c2670_wire_468,
c2670_wire_469,
c2670_wire_470,
c2670_wire_471,
c2670_wire_472,
c2670_wire_473,
c2670_wire_474,
c2670_wire_475,
c2670_wire_476,
c2670_wire_477,
c2670_wire_478,
c2670_wire_479,
c2670_wire_480,
c2670_wire_481,
c2670_wire_482,
c2670_wire_483,
c2670_wire_484,
c2670_wire_485,
c2670_wire_486,
c2670_wire_487,
c2670_wire_488,
c2670_wire_489,
c2670_wire_490,
c2670_wire_491,
c2670_wire_492,
c2670_wire_493,
c2670_wire_494,
c2670_wire_495,
c2670_wire_496,
c2670_wire_497,
c2670_wire_498,
c2670_wire_499,
c2670_wire_500,
c2670_wire_501,
c2670_wire_502,
c2670_wire_503,
c2670_wire_504,
c2670_wire_505,
c2670_wire_506,
c2670_wire_507,
c2670_wire_508,
c2670_wire_509,
c2670_wire_510,
c2670_wire_511,
c2670_wire_512,
c2670_wire_513,
c2670_wire_514,
c2670_wire_515,
c2670_wire_516,
c2670_wire_517,
c2670_wire_518,
c2670_wire_519,
c2670_wire_520,
c2670_wire_521,
c2670_wire_522,
c2670_wire_523,
c2670_wire_524,
c2670_wire_525,
c2670_wire_526,
c2670_wire_527,
c2670_wire_528,
c2670_wire_529,
c2670_wire_530,
c2670_wire_531,
c2670_wire_532,
c2670_wire_533,
c2670_wire_534,
c2670_wire_535,
c2670_wire_536,
c2670_wire_537,
c2670_wire_538,
c2670_wire_539,
c2670_wire_540,
c2670_wire_541,
c2670_wire_542,
c2670_wire_543,
c2670_wire_544,
c2670_wire_545,
c2670_wire_546,
c2670_wire_547,
c2670_wire_548,
c2670_wire_549,
c2670_wire_550,
c2670_wire_551,
c2670_wire_552,
c2670_wire_553,
c2670_wire_554,
c2670_wire_555,
c2670_wire_556,
c2670_wire_557,
c2670_wire_558,
c2670_wire_559,
c2670_wire_560,
c2670_wire_561,
c2670_wire_562,
c2670_wire_563,
c2670_wire_564,
c2670_wire_565,
c2670_wire_566,
c2670_wire_567,
c2670_wire_568,
c2670_wire_569,
c2670_wire_570,
c2670_wire_571,
c2670_wire_572,
c2670_wire_573,
c2670_wire_574,
c2670_wire_575,
c2670_wire_576,
c2670_wire_577,
c2670_wire_578,
c2670_wire_579,
c2670_wire_580,
c2670_wire_581,
c2670_wire_582,
c2670_wire_583,
c2670_wire_584,
c2670_wire_585,
c2670_wire_586,
c2670_wire_587,
c2670_wire_588,
c2670_wire_589,
c2670_wire_590,
c2670_wire_591,
c2670_wire_592,
c2670_wire_593,
c2670_wire_594,
c2670_wire_595,
c2670_wire_596,
c2670_wire_597,
c2670_wire_598,
c2670_wire_599,
c2670_wire_600,
c2670_wire_601,
c2670_wire_602,
c2670_wire_603,
c2670_wire_604,
c2670_wire_605,
c2670_wire_606,
c2670_wire_607,
c2670_wire_608,
c2670_wire_609,
c2670_wire_610,
c2670_wire_611,
c2670_wire_612,
c2670_wire_613,
c2670_wire_614,
c2670_wire_615,
c2670_wire_616,
c2670_wire_617,
c2670_wire_618,
c2670_wire_619,
c2670_wire_620,
c2670_wire_621,
c2670_wire_622,
c2670_wire_623,
c2670_wire_624,
c2670_wire_625,
c2670_wire_626,
c2670_wire_627,
c2670_wire_628,
c2670_wire_629,
c2670_wire_630,
c2670_wire_631,
c2670_wire_632,
c2670_wire_633,
c2670_wire_634,
c2670_wire_635,
c2670_wire_636,
c2670_wire_637,
c2670_wire_638,
c2670_wire_639,
c2670_wire_640,
c2670_wire_641,
c2670_wire_642,
c2670_wire_643,
c2670_wire_644,
c2670_wire_645,
c2670_wire_646,
c2670_wire_647,
c2670_wire_648,
c2670_wire_649,
c2670_wire_650,
c2670_wire_651,
c2670_wire_652,
c2670_wire_653,
c2670_wire_654,
c2670_wire_655,
c2670_wire_656,
c2670_wire_657,
c2670_wire_658,
c2670_wire_659,
c2670_wire_660,
c2670_wire_661,
c2670_wire_662,
c2670_wire_663,
c2670_wire_664,
c2670_wire_665,
c2670_wire_666,
c2670_wire_667,
c2670_wire_668,
c2670_wire_669,
c2670_wire_670,
c2670_wire_671,
c2670_wire_672,
c2670_wire_673,
c2670_wire_674,
c2670_wire_675,
c2670_wire_676,
c2670_wire_677,
c2670_wire_678,
c2670_wire_679,
c2670_wire_680,
c2670_wire_681,
c2670_wire_682,
c2670_wire_683,
c2670_wire_684,
c2670_wire_685,
c2670_wire_686,
c2670_wire_687,
c2670_wire_688,
c2670_wire_689,
c2670_wire_690,
c2670_wire_691,
c2670_wire_692,
c2670_wire_693,
c2670_wire_694,
c2670_wire_695,
c2670_wire_696,
c2670_wire_697,
c2670_wire_698,
c2670_wire_699,
c2670_wire_700,
c2670_wire_701,
c2670_wire_702,
c2670_wire_703,
c2670_wire_704,
c2670_wire_705,
c2670_wire_706,
c2670_wire_707,
c2670_wire_708,
c2670_wire_709,
c2670_wire_710,
c2670_wire_711,
c2670_wire_712,
c2670_wire_713,
c2670_wire_714,
c2670_wire_715,
c2670_wire_716,
c2670_wire_717,
c2670_wire_718,
c2670_wire_719,
c2670_wire_720,
c2670_wire_721,
c2670_wire_722,
c2670_wire_723,
c2670_wire_724,
c2670_wire_725,
c2670_wire_726,
c2670_wire_727,
c2670_wire_728,
c2670_wire_729,
c2670_wire_730,
c2670_wire_731,
c2670_wire_732,
c2670_wire_733,
c2670_wire_734,
c2670_wire_735,
c2670_wire_736,
c2670_wire_737,
c2670_wire_738,
c2670_wire_739,
c2670_wire_740,
c2670_wire_741,
c2670_wire_742,
c2670_wire_743,
c2670_wire_744,
c2670_wire_745,
c2670_wire_746,
c2670_wire_747,
c2670_wire_748,
c2670_wire_749,
c2670_wire_750,
c2670_wire_751,
c2670_wire_752,
c2670_wire_753,
c2670_wire_754,
c2670_wire_755,
c2670_wire_756,
c2670_wire_757,
c2670_wire_758,
c2670_wire_759,
c2670_wire_760,
c2670_wire_761,
c2670_wire_762,
c2670_wire_763,
c2670_wire_764,
c2670_wire_765,
c2670_wire_766,
c2670_wire_767,
c2670_wire_768,
c2670_wire_769,
c2670_wire_770,
c2670_wire_771,
c2670_wire_772,
c2670_wire_773,
c2670_wire_774,
c2670_wire_775,
c2670_wire_776,
c2670_wire_777,
c2670_wire_778,
c2670_wire_779,
c2670_wire_780,
c2670_wire_781,
c2670_wire_782,
c2670_wire_783,
c2670_wire_784,
c2670_wire_785,
c2670_wire_786,
c2670_wire_787,
c2670_wire_788,
c2670_wire_789,
c2670_wire_790,
c2670_wire_791,
c2670_wire_792,
c2670_wire_793,
c2670_wire_794,
c2670_wire_795,
c2670_wire_796,
c2670_wire_797,
c2670_wire_798,
c2670_wire_799,
c2670_wire_800,
c2670_wire_801,
c2670_wire_802,
c2670_wire_803,
c2670_wire_804,
c2670_wire_805,
c2670_wire_806,
c2670_wire_807,
c2670_wire_808,
c2670_wire_809,
c2670_wire_810,
c2670_wire_811,
c2670_wire_812,
c2670_wire_813,
c2670_wire_814,
c2670_wire_815,
c2670_wire_816,
c2670_wire_817,
c2670_wire_818,
c2670_wire_819,
c2670_wire_820,
c2670_wire_821,
c2670_wire_822,
c2670_wire_823,
c2670_wire_824,
c2670_wire_825,
c2670_wire_826,
c2670_wire_827,
c2670_wire_828,
c2670_wire_829,
c2670_wire_830,
c2670_wire_831,
c2670_wire_832,
c2670_wire_833,
c2670_wire_834,
c2670_wire_835,
c2670_wire_836,
c2670_wire_837,
c2670_wire_838,
c2670_wire_839,
c2670_wire_840,
c2670_wire_841,
c2670_wire_842,
c2670_wire_843,
c2670_wire_844,
c2670_wire_845,
c2670_wire_846,
c2670_wire_847,
c2670_wire_848,
c2670_wire_849,
c2670_wire_850,
c2670_wire_851,
c2670_wire_852,
c2670_wire_853,
c2670_wire_854,
c2670_wire_855,
c2670_wire_856,
c2670_wire_857,
c2670_wire_858,
c2670_wire_859,
c2670_wire_860,
c2670_wire_861,
c2670_wire_862,
c2670_wire_863,
c2670_wire_864,
c2670_wire_865,
c2670_wire_866,
c2670_wire_867,
c2670_wire_868,
c2670_wire_869,
c2670_wire_870,
c2670_wire_871,
c2670_wire_872,
c2670_wire_873,
c2670_wire_874,
c2670_wire_875,
c2670_wire_876,
c2670_wire_877,
c2670_wire_878,
c2670_wire_879,
c2670_wire_880,
c2670_wire_881,
c2670_wire_882,
c2670_wire_883,
c2670_wire_884,
c2670_wire_885,
c2670_wire_886,
c2670_wire_887,
c2670_wire_888,
c2670_wire_889,
c2670_wire_890,
c2670_wire_891,
c2670_wire_892,
c2670_wire_893,
c2670_wire_894,
c2670_wire_895,
c2670_wire_896,
c2670_wire_897,
c2670_wire_898,
c2670_wire_899,
c2670_wire_900,
c2670_wire_901,
c2670_wire_902,
c2670_wire_903,
c2670_wire_904,
c2670_wire_905,
c2670_wire_906,
c2670_wire_907,
c2670_wire_908,
c2670_wire_909,
c2670_wire_910,
c2670_wire_911,
c2670_wire_912,
c2670_wire_913,
c2670_wire_914,
c2670_wire_915,
c2670_wire_916,
c2670_wire_917,
c2670_wire_918,
c2670_wire_919,
c2670_wire_920,
c2670_wire_921,
c2670_wire_922,
c2670_wire_923,
c2670_wire_924,
c2670_wire_925,
c2670_wire_926,
c2670_wire_927,
c2670_wire_928,
c2670_wire_929,
c2670_wire_930,
c2670_wire_931,
c2670_wire_932,
c2670_wire_933,
c2670_wire_934,
c2670_wire_935,
c2670_wire_936,
c2670_wire_937,
c2670_wire_938,
c2670_wire_939,
c2670_wire_940,
c2670_wire_941,
c2670_wire_942,
c2670_wire_943,
c2670_wire_944,
c2670_wire_945,
c2670_wire_946,
c2670_wire_947,
c2670_wire_948,
c2670_wire_949,
c2670_wire_950,
c2670_wire_951,
c2670_wire_952,
c2670_wire_953,
c2670_wire_954,
c2670_wire_955,
c2670_wire_956,
c2670_wire_957,
c2670_wire_958,
c2670_wire_959,
c2670_wire_960,
c2670_wire_961,
c2670_wire_962,
c2670_wire_963,
c2670_wire_964,
c2670_wire_965,
c2670_wire_966,
c2670_wire_967,
c2670_wire_968,
c2670_wire_969,
c2670_wire_970,
c2670_wire_971,
c2670_wire_972,
c2670_wire_973,
c2670_wire_974,
c2670_wire_975,
c2670_wire_976,
c2670_wire_977,
c2670_wire_978,
c2670_wire_979,
c2670_wire_980,
c2670_wire_981,
c2670_wire_982,
c2670_wire_5_0,
c2670_wire_5_1,
c2670_wire_5_2,
c2670_wire_5_3,
c2670_wire_5_4,
c2670_wire_5_5,
c2670_wire_5_6,
c2670_wire_5_7,
c2670_wire_5_8,
c2670_wire_34_0,
c2670_wire_34_1,
c2670_wire_34_2,
c2670_wire_34_3,
c2670_wire_35_0,
c2670_wire_35_1,
c2670_wire_35_2,
c2670_wire_35_3,
c2670_wire_35_4,
c2670_wire_35_5,
c2670_wire_35_6,
c2670_wire_35_7,
c2670_wire_35_8,
c2670_wire_35_9,
c2670_wire_35_10,
c2670_wire_35_11,
c2670_wire_36_0,
c2670_wire_36_1,
c2670_wire_36_2,
c2670_wire_36_3,
c2670_wire_36_4,
c2670_wire_36_5,
c2670_wire_36_6,
c2670_wire_36_7,
c2670_wire_36_8,
c2670_wire_36_9,
c2670_wire_36_10,
c2670_wire_91_0,
c2670_wire_91_1,
c2670_wire_91_2,
c2670_wire_91_3,
c2670_wire_91_4,
c2670_wire_91_5,
c2670_wire_91_6,
c2670_wire_91_7,
c2670_wire_91_8,
c2670_wire_91_9,
c2670_wire_110_0,
c2670_wire_110_1,
c2670_wire_110_2,
c2670_wire_110_3,
c2670_wire_110_4,
c2670_wire_110_5,
c2670_wire_110_6,
c2670_wire_126_0,
c2670_wire_126_1,
c2670_wire_126_2,
c2670_wire_126_3,
c2670_wire_126_4,
c2670_wire_126_5,
c2670_wire_126_6,
c2670_wire_126_7,
c2670_wire_126_8,
c2670_wire_147_0,
c2670_wire_147_1,
c2670_wire_147_2,
c2670_wire_147_3,
c2670_wire_147_4,
c2670_wire_147_5,
c2670_wire_147_6,
c2670_wire_147_7,
c2670_wire_157_0,
c2670_wire_157_1,
c2670_wire_157_2,
c2670_wire_157_3,
c2670_wire_157_4,
c2670_wire_173_0,
c2670_wire_173_1,
c2670_wire_173_2,
c2670_wire_173_3,
c2670_wire_173_4,
c2670_wire_173_5,
c2670_wire_173_6,
c2670_wire_173_7,
c2670_wire_181_0,
c2670_wire_181_1,
c2670_wire_181_2,
c2670_wire_181_3,
c2670_wire_181_4,
c2670_wire_181_5,
c2670_wire_181_6,
c2670_wire_209_0,
c2670_wire_209_1,
c2670_wire_209_2,
c2670_wire_209_3,
c2670_wire_209_4,
c2670_wire_209_5,
c2670_wire_209_6,
c2670_wire_211_0,
c2670_wire_211_1,
c2670_wire_211_2,
c2670_wire_211_3,
c2670_wire_211_4,
c2670_wire_251_0,
c2670_wire_251_1,
c2670_wire_251_2,
c2670_wire_251_3,
c2670_wire_251_4,
c2670_wire_275_0,
c2670_wire_275_1,
c2670_wire_276_0,
c2670_wire_276_1,
c2670_wire_277_0,
c2670_wire_277_1,
c2670_wire_277_2,
c2670_wire_277_3,
c2670_wire_277_4,
c2670_wire_277_5,
c2670_wire_297_0,
c2670_wire_297_1,
c2670_wire_297_2,
c2670_wire_297_3,
c2670_wire_297_4,
c2670_wire_297_5,
c2670_wire_297_6,
c2670_wire_297_7,
c2670_wire_318_0,
c2670_wire_318_1,
c2670_wire_298_0,
c2670_wire_298_1,
c2670_wire_298_2,
c2670_wire_298_3,
c2670_wire_298_4,
c2670_wire_298_5,
c2670_wire_298_6,
c2670_wire_183_0,
c2670_wire_183_1,
c2670_wire_183_2,
c2670_wire_183_3,
c2670_wire_370_0,
c2670_wire_370_1,
c2670_wire_375_0,
c2670_wire_375_1,
c2670_wire_378_0,
c2670_wire_378_1,
c2670_wire_382_0,
c2670_wire_382_1,
c2670_wire_386_0,
c2670_wire_386_1,
c2670_wire_389_0,
c2670_wire_389_1,
c2670_wire_392_0,
c2670_wire_392_1,
c2670_wire_396_0,
c2670_wire_396_1,
c2670_wire_401_0,
c2670_wire_401_1,
c2670_wire_406_0,
c2670_wire_406_1,
c2670_wire_406_2,
c2670_wire_406_3,
c2670_wire_428_0,
c2670_wire_428_1,
c2670_wire_428_2,
c2670_wire_416_0,
c2670_wire_416_1,
c2670_wire_24_0,
c2670_wire_24_1,
c2670_wire_24_2,
c2670_wire_24_3,
c2670_wire_24_4,
c2670_wire_24_5,
c2670_wire_24_6,
c2670_wire_24_7,
c2670_wire_24_8,
c2670_wire_24_9,
c2670_wire_24_10,
c2670_wire_24_11,
c2670_wire_24_12,
c2670_wire_24_13,
c2670_wire_24_14,
c2670_wire_24_15,
c2670_wire_24_16,
c2670_wire_24_17,
c2670_wire_24_18,
c2670_wire_24_19,
c2670_wire_13_0,
c2670_wire_13_1,
c2670_wire_13_2,
c2670_wire_13_3,
c2670_wire_13_4,
c2670_wire_13_5,
c2670_wire_434_0,
c2670_wire_434_1,
c2670_wire_441_0,
c2670_wire_441_1,
c2670_wire_441_2,
c2670_wire_441_3,
c2670_wire_441_4,
c2670_wire_441_5,
c2670_wire_441_6,
c2670_wire_441_7,
c2670_wire_441_8,
c2670_wire_441_9,
c2670_wire_441_10,
c2670_wire_441_11,
c2670_wire_441_12,
c2670_wire_441_13,
c2670_wire_441_14,
c2670_wire_441_15,
c2670_wire_441_16,
c2670_wire_441_17,
c2670_wire_441_18,
c2670_wire_441_19,
c2670_wire_441_20,
c2670_wire_441_21,
c2670_wire_441_22,
c2670_wire_441_23,
c2670_wire_441_24,
c2670_wire_441_25,
c2670_wire_441_26,
c2670_wire_441_27,
c2670_wire_20_0,
c2670_wire_20_1,
c2670_wire_20_2,
c2670_wire_20_3,
c2670_wire_20_4,
c2670_wire_20_5,
c2670_wire_20_6,
c2670_wire_20_7,
c2670_wire_20_8,
c2670_wire_20_9,
c2670_wire_20_10,
c2670_wire_20_11,
c2670_wire_20_12,
c2670_wire_20_13,
c2670_wire_20_14,
c2670_wire_20_15,
c2670_wire_20_16,
c2670_wire_20_17,
c2670_wire_20_18,
c2670_wire_20_19,
c2670_wire_20_20,
c2670_wire_20_21,
c2670_wire_20_22,
c2670_wire_20_23,
c2670_wire_20_24,
c2670_wire_20_25,
c2670_wire_20_26,
c2670_wire_20_27,
c2670_wire_20_28,
c2670_wire_20_29,
c2670_wire_20_30,
c2670_wire_20_31,
c2670_wire_20_32,
c2670_wire_20_33,
c2670_wire_20_34,
c2670_wire_20_35,
c2670_wire_20_36,
c2670_wire_20_37,
c2670_wire_20_38,
c2670_wire_419_0,
c2670_wire_419_1,
c2670_wire_419_2,
c2670_wire_419_3,
c2670_wire_419_4,
c2670_wire_419_5,
c2670_wire_450_0,
c2670_wire_450_1,
c2670_wire_450_2,
c2670_wire_450_3,
c2670_wire_453_0,
c2670_wire_453_1,
c2670_wire_453_2,
c2670_wire_453_3,
c2670_wire_453_4,
c2670_wire_453_5,
c2670_wire_453_6,
c2670_wire_453_7,
c2670_wire_464_0,
c2670_wire_464_1,
c2670_wire_465_0,
c2670_wire_465_1,
c2670_wire_465_2,
c2670_wire_465_3,
c2670_wire_465_4,
c2670_wire_466_0,
c2670_wire_466_1,
c2670_wire_466_2,
c2670_wire_466_3,
c2670_wire_466_4,
c2670_wire_471_0,
c2670_wire_471_1,
c2670_wire_371_0,
c2670_wire_371_1,
c2670_wire_371_2,
c2670_wire_371_3,
c2670_wire_371_4,
c2670_wire_371_5,
c2670_wire_473_0,
c2670_wire_473_1,
c2670_wire_483_0,
c2670_wire_483_1,
c2670_wire_483_2,
c2670_wire_483_3,
c2670_wire_483_4,
c2670_wire_484_0,
c2670_wire_484_1,
c2670_wire_497_0,
c2670_wire_497_1,
c2670_wire_489_0,
c2670_wire_489_1,
c2670_wire_489_2,
c2670_wire_489_3,
c2670_wire_489_4,
c2670_wire_489_5,
c2670_wire_489_6,
c2670_wire_525_0,
c2670_wire_525_1,
c2670_wire_525_2,
c2670_wire_525_3,
c2670_wire_525_4,
c2670_wire_526_0,
c2670_wire_526_1,
c2670_wire_526_2,
c2670_wire_526_3,
c2670_wire_526_4,
c2670_wire_526_5,
c2670_wire_526_6,
c2670_wire_526_7,
c2670_wire_526_8,
c2670_wire_526_9,
c2670_wire_526_10,
c2670_wire_526_11,
c2670_wire_526_12,
c2670_wire_526_13,
c2670_wire_526_14,
c2670_wire_526_15,
c2670_wire_526_16,
c2670_wire_526_17,
c2670_wire_526_18,
c2670_wire_526_19,
c2670_wire_526_20,
c2670_wire_526_21,
c2670_wire_526_22,
c2670_wire_526_23,
c2670_wire_552_0,
c2670_wire_552_1,
c2670_wire_552_2,
c2670_wire_552_3,
c2670_wire_552_4,
c2670_wire_552_5,
c2670_wire_552_6,
c2670_wire_459_0,
c2670_wire_459_1,
c2670_wire_459_2,
c2670_wire_477_0,
c2670_wire_477_1,
c2670_wire_477_2,
c2670_wire_477_3,
c2670_wire_477_4,
c2670_wire_477_5,
c2670_wire_477_6,
c2670_wire_557_0,
c2670_wire_557_1,
c2670_wire_557_2,
c2670_wire_557_3,
c2670_wire_557_4,
c2670_wire_557_5,
c2670_wire_557_6,
c2670_wire_284_0,
c2670_wire_284_1,
c2670_wire_284_2,
c2670_wire_284_3,
c2670_wire_284_4,
c2670_wire_284_5,
c2670_wire_284_6,
c2670_wire_284_7,
c2670_wire_302_0,
c2670_wire_302_1,
c2670_wire_302_2,
c2670_wire_302_3,
c2670_wire_302_4,
c2670_wire_302_5,
c2670_wire_302_6,
c2670_wire_302_7,
c2670_wire_302_8,
c2670_wire_8_0,
c2670_wire_8_1,
c2670_wire_8_2,
c2670_wire_8_3,
c2670_wire_8_4,
c2670_wire_571_0,
c2670_wire_571_1,
c2670_wire_571_2,
c2670_wire_329_0,
c2670_wire_329_1,
c2670_wire_329_2,
c2670_wire_329_3,
c2670_wire_329_4,
c2670_wire_329_5,
c2670_wire_329_6,
c2670_wire_347_0,
c2670_wire_347_1,
c2670_wire_347_2,
c2670_wire_347_3,
c2670_wire_347_4,
c2670_wire_347_5,
c2670_wire_347_6,
c2670_wire_347_7,
c2670_wire_481_0,
c2670_wire_481_1,
c2670_wire_574_0,
c2670_wire_574_1,
c2670_wire_574_2,
c2670_wire_574_3,
c2670_wire_574_4,
c2670_wire_574_5,
c2670_wire_585_0,
c2670_wire_585_1,
c2670_wire_585_2,
c2670_wire_585_3,
c2670_wire_586_0,
c2670_wire_586_1,
c2670_wire_586_2,
c2670_wire_586_3,
c2670_wire_586_4,
c2670_wire_586_5,
c2670_wire_586_6,
c2670_wire_587_0,
c2670_wire_587_1,
c2670_wire_593_0,
c2670_wire_593_1,
c2670_wire_593_2,
c2670_wire_594_0,
c2670_wire_594_1,
c2670_wire_594_2,
c2670_wire_596_0,
c2670_wire_596_1,
c2670_wire_596_2,
c2670_wire_596_3,
c2670_wire_597_0,
c2670_wire_597_1,
c2670_wire_597_2,
c2670_wire_597_3,
c2670_wire_597_4,
c2670_wire_216_0,
c2670_wire_216_1,
c2670_wire_216_2,
c2670_wire_216_3,
c2670_wire_216_4,
c2670_wire_216_5,
c2670_wire_216_6,
c2670_wire_216_7,
c2670_wire_234_0,
c2670_wire_234_1,
c2670_wire_234_2,
c2670_wire_234_3,
c2670_wire_234_4,
c2670_wire_234_5,
c2670_wire_234_6,
c2670_wire_234_7,
c2670_wire_255_0,
c2670_wire_255_1,
c2670_wire_255_2,
c2670_wire_255_3,
c2670_wire_607_0,
c2670_wire_607_1,
c2670_wire_607_2,
c2670_wire_607_3,
c2670_wire_607_4,
c2670_wire_197_0,
c2670_wire_197_1,
c2670_wire_197_2,
c2670_wire_197_3,
c2670_wire_197_4,
c2670_wire_197_5,
c2670_wire_197_6,
c2670_wire_197_7,
c2670_wire_197_8,
c2670_wire_197_9,
c2670_wire_197_10,
c2670_wire_197_11,
c2670_wire_197_12,
c2670_wire_197_13,
c2670_wire_197_14,
c2670_wire_197_15,
c2670_wire_197_16,
c2670_wire_197_17,
c2670_wire_195_0,
c2670_wire_195_1,
c2670_wire_195_2,
c2670_wire_195_3,
c2670_wire_195_4,
c2670_wire_195_5,
c2670_wire_195_6,
c2670_wire_195_7,
c2670_wire_195_8,
c2670_wire_195_9,
c2670_wire_195_10,
c2670_wire_195_11,
c2670_wire_195_12,
c2670_wire_195_13,
c2670_wire_195_14,
c2670_wire_195_15,
c2670_wire_195_16,
c2670_wire_195_17,
c2670_wire_195_18,
c2670_wire_195_19,
c2670_wire_195_20,
c2670_wire_195_21,
c2670_wire_195_22,
c2670_wire_195_23,
c2670_wire_195_24,
c2670_wire_195_25,
c2670_wire_195_26,
c2670_wire_195_27,
c2670_wire_195_28,
c2670_wire_195_29,
c2670_wire_195_30,
c2670_wire_195_31,
c2670_wire_195_32,
c2670_wire_195_33,
c2670_wire_195_34,
c2670_wire_195_35,
c2670_wire_449_0,
c2670_wire_449_1,
c2670_wire_614_0,
c2670_wire_614_1,
c2670_wire_616_0,
c2670_wire_616_1,
c2670_wire_523_0,
c2670_wire_523_1,
c2670_wire_617_0,
c2670_wire_617_1,
c2670_wire_622_0,
c2670_wire_622_1,
c2670_wire_623_0,
c2670_wire_623_1,
c2670_wire_624_0,
c2670_wire_624_1,
c2670_wire_626_0,
c2670_wire_626_1,
c2670_wire_629_0,
c2670_wire_629_1,
c2670_wire_630_0,
c2670_wire_630_1,
c2670_wire_632_0,
c2670_wire_632_1,
c2670_wire_410_0,
c2670_wire_410_1,
c2670_wire_410_2,
c2670_wire_410_3,
c2670_wire_634_0,
c2670_wire_634_1,
c2670_wire_634_2,
c2670_wire_634_3,
c2670_wire_610_0,
c2670_wire_610_1,
c2670_wire_610_2,
c2670_wire_610_3,
c2670_wire_505_0,
c2670_wire_505_1,
c2670_wire_513_0,
c2670_wire_513_1,
c2670_wire_716_0,
c2670_wire_716_1,
c2670_wire_716_2,
c2670_wire_716_3,
c2670_wire_719_0,
c2670_wire_719_1,
c2670_wire_518_0,
c2670_wire_518_1,
c2670_wire_732_0,
c2670_wire_732_1,
c2670_wire_742_0,
c2670_wire_742_1,
c2670_wire_744_0,
c2670_wire_744_1,
c2670_wire_755_0,
c2670_wire_755_1,
c2670_wire_755_2,
c2670_wire_758_0,
c2670_wire_758_1,
c2670_wire_762_0,
c2670_wire_762_1,
c2670_wire_762_2,
c2670_wire_764_0,
c2670_wire_764_1,
c2670_wire_769_0,
c2670_wire_769_1,
c2670_wire_771_0,
c2670_wire_771_1,
c2670_wire_452_0,
c2670_wire_452_1,
c2670_wire_670_0,
c2670_wire_670_1,
c2670_wire_693_0,
c2670_wire_693_1,
c2670_wire_693_2,
c2670_wire_693_3,
c2670_wire_676_0,
c2670_wire_676_1,
c2670_wire_779_0,
c2670_wire_779_1,
c2670_wire_779_2,
c2670_wire_779_3,
c2670_wire_787_0,
c2670_wire_787_1,
c2670_wire_787_2,
c2670_wire_787_3,
c2670_wire_792_0,
c2670_wire_792_1,
c2670_wire_792_2,
c2670_wire_792_3,
c2670_wire_796_0,
c2670_wire_796_1,
c2670_wire_805_0,
c2670_wire_805_1,
c2670_wire_805_2,
c2670_wire_805_3,
c2670_wire_782_0,
c2670_wire_782_1,
c2670_wire_782_2,
c2670_wire_782_3,
c2670_wire_759_0,
c2670_wire_759_1,
c2670_wire_759_2,
c2670_wire_765_0,
c2670_wire_765_1,
c2670_wire_765_2,
c2670_wire_806_0,
c2670_wire_806_1,
c2670_wire_488_0,
c2670_wire_488_1,
c2670_wire_488_2,
c2670_wire_488_3,
c2670_wire_488_4,
c2670_wire_488_5,
c2670_wire_488_6,
c2670_wire_488_7,
c2670_wire_488_8,
c2670_wire_488_9,
c2670_wire_488_10,
c2670_wire_488_11,
c2670_wire_488_12,
c2670_wire_488_13,
c2670_wire_488_14,
c2670_wire_488_15,
c2670_wire_488_16,
c2670_wire_488_17,
c2670_wire_827_0,
c2670_wire_827_1,
c2670_wire_846_0,
c2670_wire_846_1,
c2670_wire_846_2,
c2670_wire_846_3,
c2670_wire_850_0,
c2670_wire_850_1,
c2670_wire_664_0,
c2670_wire_664_1,
c2670_wire_854_0,
c2670_wire_854_1,
c2670_wire_858_0,
c2670_wire_858_1,
c2670_wire_862_0,
c2670_wire_862_1,
c2670_wire_879_0,
c2670_wire_879_1,
c2670_wire_864_0,
c2670_wire_864_1,
c2670_wire_577_0,
c2670_wire_577_1,
c2670_wire_899_0,
c2670_wire_899_1,
c2670_wire_899_2,
c2670_wire_928_0,
c2670_wire_928_1,
c2670_wire_929_0,
c2670_wire_929_1,
c2670_wire_934_0,
c2670_wire_934_1,
c2670_wire_934_2,
c2670_wire_954_0,
c2670_wire_954_1,
c2670_wire_961_0,
c2670_wire_961_1,
c2670_wire_963_0,
c2670_wire_963_1,
c2670_wire_964_0,
c2670_wire_964_1,
c2670_wire_970_0,
c2670_wire_970_1,
c2670_wire_602_0,
c2670_wire_602_1,
c2670_wire_604_0,
c2670_wire_604_1,
c2670_wire_835_0,
c2670_wire_835_1,
c2670_wire_187_0,
c2670_wire_187_1,
c2670_wire_319_0,
c2670_wire_319_1,
c2670_wire_955_0,
c2670_wire_955_1,
c2670_wire_510_0,
c2670_wire_510_1,
c2670_wire_943_0,
c2670_wire_943_1,
c2670_wire_500_0,
c2670_wire_500_1,
c2670_wire_939_0,
c2670_wire_939_1,
c2670_wire_320_0,
c2670_wire_320_1,
c2670_wire_582_0,
c2670_wire_582_1,
c2670_wire_579_0,
c2670_wire_579_1,
c2670_wire_580_0,
c2670_wire_580_1,
c2670_wire_438_0,
c2670_wire_438_1,
c2670_wire_438_2,
c2670_wire_321_0,
c2670_wire_321_1,
c2670_wire_619_0,
c2670_wire_619_1,
c2670_wire_619_2,
c2670_wire_619_3,
c2670_wire_757_0,
c2670_wire_757_1,
c2670_wire_757_2,
c2670_wire_757_3,
c2670_wire_757_4,
c2670_wire_757_5,
c2670_wire_757_6,
c2670_wire_757_7,
c2670_wire_945_0,
c2670_wire_945_1,
c2670_wire_941_0,
c2670_wire_941_1,
c2670_wire_420_0,
c2670_wire_420_1,
c2670_wire_420_2,
c2670_wire_420_3,
G1_net_0,
G2_net_0,
G3_net_0,
G4_net_0,
G5_net_0,
G6_net_0,
G7_net_0,
G8_net_0,
G9_net_0,
G10_net_0,
G11_net_0,
G12_net_0,
G13_net_0,
G14_net_0,
G15_net_0,
G16_net_0,
G17_net_0,
G18_net_0,
G19_net_0,
G20_net_0,
G21_net_0,
G22_net_0,
G23_net_0,
G24_net_0,
G25_net_0,
G26_net_0,
G27_net_0,
G28_net_0,
G29_net_0,
G30_net_0,
G31_net_0,
G32_net_0,
G33_net_0,
G34_net_0,
G35_net_0,
G36_net_0,
G37_net_0,
G38_net_0,
G39_net_0,
G40_net_0,
G41_net_0,
G42_net_0,
G43_net_0,
G44_net_0,
G45_net_0,
G46_net_0,
G47_net_0,
G48_net_0,
G49_net_0,
G50_net_0,
G51_net_0,
G52_net_0,
G53_net_0,
G54_net_0,
G55_net_0,
G56_net_0,
G57_net_0,
G58_net_0,
G59_net_0,
G60_net_0,
G61_net_0,
G62_net_0,
G63_net_0,
G64_net_0,
G65_net_0,
G66_net_0,
G67_net_0,
G68_net_0,
G69_net_0,
G70_net_0,
G71_net_0,
G72_net_0,
G73_net_0,
G74_net_0,
G75_net_0,
G76_net_0,
G77_net_0,
G78_net_0,
G79_net_0,
G80_net_0,
G81_net_0,
G82_net_0,
G83_net_0,
G84_net_0,
G85_net_0,
G86_net_0,
G87_net_0,
G88_net_0,
G89_net_0,
G90_net_0,
G91_net_0,
G92_net_0,
G93_net_0,
G94_net_0,
G95_net_0,
G96_net_0,
G97_net_0,
G98_net_0,
G99_net_0,
G100_net_0,
G101_net_0,
G102_net_0,
G103_net_0,
G104_net_0,
G105_net_0,
G106_net_0,
G107_net_0,
G108_net_0,
G109_net_0,
G110_net_0,
G111_net_0,
G112_net_0,
G113_net_0,
G114_net_0,
G115_net_0,
G116_net_0,
G117_net_0,
G118_net_0,
G119_net_0,
G120_net_0,
G121_net_0,
G122_net_0,
G123_net_0,
G124_net_0,
G125_net_0,
G126_net_0,
G127_net_0,
G128_net_0,
G129_net_0,
G130_net_0,
G131_net_0,
G132_net_0,
G133_net_0,
G134_net_0,
G135_net_0,
G136_net_0,
G137_net_0,
G138_net_0,
G139_net_0,
G140_net_0,
G141_net_0,
G142_net_0,
G143_net_0,
G144_net_0,
G145_net_0,
G146_net_0,
G147_net_0,
G148_net_0,
G149_net_0,
G150_net_0,
G151_net_0,
G152_net_0,
G153_net_0,
G154_net_0,
G155_net_0,
G156_net_0,
G157_net_0,
G2531_net_0,
G2532_net_0,
G2533_net_0,
G2534_net_0,
G2535_net_0,
G2536_net_0,
G2537_net_0,
G2538_net_0,
G2539_net_0,
G2540_net_0,
G2541_net_0,
G2542_net_0,
G2543_net_0,
G2544_net_0,
G2545_net_0,
G2546_net_0,
G2547_net_0,
G2548_net_0,
G2549_net_0,
G2550_net_0,
G2551_net_0,
G2552_net_0,
G2553_net_0,
G2554_net_0,
G2555_net_0,
G2556_net_0,
G2557_net_0,
G2558_net_0,
G2559_net_0,
G2560_net_0,
G2561_net_0,
G2562_net_0,
G2563_net_0,
G2564_net_0,
G2565_net_0,
G2566_net_0,
G2567_net_0,
G2568_net_0,
G2569_net_0,
G2570_net_0,
G2571_net_0,
G2572_net_0,
G2573_net_0,
G2574_net_0,
G2575_net_0,
G2576_net_0,
G2577_net_0,
G2578_net_0,
G2579_net_0,
G2580_net_0,
G2581_net_0,
G2582_net_0,
G2583_net_0,
G2584_net_0,
G2585_net_0,
G2586_net_0,
G2587_net_0,
G2588_net_0,
G2589_net_0,
G2590_net_0,
G2591_net_0,
G2592_net_0,
G2593_net_0,
G2594_net_0;

pin #(157) pin_0 ({G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157}, {G1_net_0, G2_net_0, G3_net_0, G4_net_0, G5_net_0, G6_net_0, G7_net_0, G8_net_0, G9_net_0, G10_net_0, G11_net_0, G12_net_0, G13_net_0, G14_net_0, G15_net_0, G16_net_0, G17_net_0, G18_net_0, G19_net_0, G20_net_0, G21_net_0, G22_net_0, G23_net_0, G24_net_0, G25_net_0, G26_net_0, G27_net_0, G28_net_0, G29_net_0, G30_net_0, G31_net_0, G32_net_0, G33_net_0, G34_net_0, G35_net_0, G36_net_0, G37_net_0, G38_net_0, G39_net_0, G40_net_0, G41_net_0, G42_net_0, G43_net_0, G44_net_0, G45_net_0, G46_net_0, G47_net_0, G48_net_0, G49_net_0, G50_net_0, G51_net_0, G52_net_0, G53_net_0, G54_net_0, G55_net_0, G56_net_0, G57_net_0, G58_net_0, G59_net_0, G60_net_0, G61_net_0, G62_net_0, G63_net_0, G64_net_0, G65_net_0, G66_net_0, G67_net_0, G68_net_0, G69_net_0, G70_net_0, G71_net_0, G72_net_0, G73_net_0, G74_net_0, G75_net_0, G76_net_0, G77_net_0, G78_net_0, G79_net_0, G80_net_0, G81_net_0, G82_net_0, G83_net_0, G84_net_0, G85_net_0, G86_net_0, G87_net_0, G88_net_0, G89_net_0, G90_net_0, G91_net_0, G92_net_0, G93_net_0, G94_net_0, G95_net_0, G96_net_0, G97_net_0, G98_net_0, G99_net_0, G100_net_0, G101_net_0, G102_net_0, G103_net_0, G104_net_0, G105_net_0, G106_net_0, G107_net_0, G108_net_0, G109_net_0, G110_net_0, G111_net_0, G112_net_0, G113_net_0, G114_net_0, G115_net_0, G116_net_0, G117_net_0, G118_net_0, G119_net_0, G120_net_0, G121_net_0, G122_net_0, G123_net_0, G124_net_0, G125_net_0, G126_net_0, G127_net_0, G128_net_0, G129_net_0, G130_net_0, G131_net_0, G132_net_0, G133_net_0, G134_net_0, G135_net_0, G136_net_0, G137_net_0, G138_net_0, G139_net_0, G140_net_0, G141_net_0, G142_net_0, G143_net_0, G144_net_0, G145_net_0, G146_net_0, G147_net_0, G148_net_0, G149_net_0, G150_net_0, G151_net_0, G152_net_0, G153_net_0, G154_net_0, G155_net_0, G156_net_0, G157_net_0});

pout #(64) pout_0 ({G2531_net_0, G2532_net_0, G2533_net_0, G2534_net_0, G2535_net_0, G2536_net_0, G2537_net_0, G2538_net_0, G2539_net_0, G2540_net_0, G2541_net_0, G2542_net_0, G2543_net_0, G2544_net_0, G2545_net_0, G2546_net_0, G2547_net_0, G2548_net_0, G2549_net_0, G2550_net_0, G2551_net_0, G2552_net_0, G2553_net_0, G2554_net_0, G2555_net_0, G2556_net_0, G2557_net_0, G2558_net_0, G2559_net_0, G2560_net_0, G2561_net_0, G2562_net_0, G2563_net_0, G2564_net_0, G2565_net_0, G2566_net_0, G2567_net_0, G2568_net_0, G2569_net_0, G2570_net_0, G2571_net_0, G2572_net_0, G2573_net_0, G2574_net_0, G2575_net_0, G2576_net_0, G2577_net_0, G2578_net_0, G2579_net_0, G2580_net_0, G2581_net_0, G2582_net_0, G2583_net_0, G2584_net_0, G2585_net_0, G2586_net_0, G2587_net_0, G2588_net_0, G2589_net_0, G2590_net_0, G2591_net_0, G2592_net_0, G2593_net_0, G2594_net_0}, {G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594});

fanout_n #(9, 0, 0) FANOUT_1 (c2670_wire_5, {c2670_wire_5_0, c2670_wire_5_1, c2670_wire_5_2, c2670_wire_5_3, c2670_wire_5_4, c2670_wire_5_5, c2670_wire_5_6, c2670_wire_5_7, c2670_wire_5_8});
fanout_n #(4, 0, 0) FANOUT_2 (c2670_wire_34, {c2670_wire_34_0, c2670_wire_34_1, c2670_wire_34_2, c2670_wire_34_3});
fanout_n #(12, 0, 0) FANOUT_3 (c2670_wire_35, {c2670_wire_35_0, c2670_wire_35_1, c2670_wire_35_2, c2670_wire_35_3, c2670_wire_35_4, c2670_wire_35_5, c2670_wire_35_6, c2670_wire_35_7, c2670_wire_35_8, c2670_wire_35_9, c2670_wire_35_10, c2670_wire_35_11});
fanout_n #(11, 0, 0) FANOUT_4 (c2670_wire_36, {c2670_wire_36_0, c2670_wire_36_1, c2670_wire_36_2, c2670_wire_36_3, c2670_wire_36_4, c2670_wire_36_5, c2670_wire_36_6, c2670_wire_36_7, c2670_wire_36_8, c2670_wire_36_9, c2670_wire_36_10});
fanout_n #(10, 0, 0) FANOUT_5 (c2670_wire_91, {c2670_wire_91_0, c2670_wire_91_1, c2670_wire_91_2, c2670_wire_91_3, c2670_wire_91_4, c2670_wire_91_5, c2670_wire_91_6, c2670_wire_91_7, c2670_wire_91_8, c2670_wire_91_9});
fanout_n #(7, 0, 0) FANOUT_6 (c2670_wire_110, {c2670_wire_110_0, c2670_wire_110_1, c2670_wire_110_2, c2670_wire_110_3, c2670_wire_110_4, c2670_wire_110_5, c2670_wire_110_6});
fanout_n #(9, 0, 0) FANOUT_7 (c2670_wire_126, {c2670_wire_126_0, c2670_wire_126_1, c2670_wire_126_2, c2670_wire_126_3, c2670_wire_126_4, c2670_wire_126_5, c2670_wire_126_6, c2670_wire_126_7, c2670_wire_126_8});
fanout_n #(8, 0, 0) FANOUT_8 (c2670_wire_147, {c2670_wire_147_0, c2670_wire_147_1, c2670_wire_147_2, c2670_wire_147_3, c2670_wire_147_4, c2670_wire_147_5, c2670_wire_147_6, c2670_wire_147_7});
fanout_n #(5, 0, 0) FANOUT_9 (c2670_wire_157, {c2670_wire_157_0, c2670_wire_157_1, c2670_wire_157_2, c2670_wire_157_3, c2670_wire_157_4});
fanout_n #(8, 0, 0) FANOUT_10 (c2670_wire_173, {c2670_wire_173_0, c2670_wire_173_1, c2670_wire_173_2, c2670_wire_173_3, c2670_wire_173_4, c2670_wire_173_5, c2670_wire_173_6, c2670_wire_173_7});
fanout_n #(7, 0, 0) FANOUT_11 (c2670_wire_181, {c2670_wire_181_0, c2670_wire_181_1, c2670_wire_181_2, c2670_wire_181_3, c2670_wire_181_4, c2670_wire_181_5, c2670_wire_181_6});
fanout_n #(7, 0, 0) FANOUT_12 (c2670_wire_209, {c2670_wire_209_0, c2670_wire_209_1, c2670_wire_209_2, c2670_wire_209_3, c2670_wire_209_4, c2670_wire_209_5, c2670_wire_209_6});
fanout_n #(5, 0, 0) FANOUT_13 (c2670_wire_211, {c2670_wire_211_0, c2670_wire_211_1, c2670_wire_211_2, c2670_wire_211_3, c2670_wire_211_4});
fanout_n #(5, 0, 0) FANOUT_14 (c2670_wire_251, {c2670_wire_251_0, c2670_wire_251_1, c2670_wire_251_2, c2670_wire_251_3, c2670_wire_251_4});
fanout_n #(2, 0, 0) FANOUT_15 (c2670_wire_275, {c2670_wire_275_0, c2670_wire_275_1});
fanout_n #(2, 0, 0) FANOUT_16 (c2670_wire_276, {c2670_wire_276_0, c2670_wire_276_1});
fanout_n #(6, 0, 0) FANOUT_17 (c2670_wire_277, {c2670_wire_277_0, c2670_wire_277_1, c2670_wire_277_2, c2670_wire_277_3, c2670_wire_277_4, c2670_wire_277_5});
fanout_n #(8, 0, 0) FANOUT_18 (c2670_wire_297, {c2670_wire_297_0, c2670_wire_297_1, c2670_wire_297_2, c2670_wire_297_3, c2670_wire_297_4, c2670_wire_297_5, c2670_wire_297_6, c2670_wire_297_7});
fanout_n #(2, 0, 0) FANOUT_19 (c2670_wire_318, {c2670_wire_318_0, c2670_wire_318_1});
fanout_n #(7, 0, 0) FANOUT_20 (c2670_wire_298, {c2670_wire_298_0, c2670_wire_298_1, c2670_wire_298_2, c2670_wire_298_3, c2670_wire_298_4, c2670_wire_298_5, c2670_wire_298_6});
fanout_n #(4, 0, 0) FANOUT_21 (c2670_wire_183, {c2670_wire_183_0, c2670_wire_183_1, c2670_wire_183_2, c2670_wire_183_3});
fanout_n #(2, 0, 0) FANOUT_22 (c2670_wire_370, {c2670_wire_370_0, c2670_wire_370_1});
fanout_n #(2, 0, 0) FANOUT_23 (c2670_wire_375, {c2670_wire_375_0, c2670_wire_375_1});
fanout_n #(2, 0, 0) FANOUT_24 (c2670_wire_378, {c2670_wire_378_0, c2670_wire_378_1});
fanout_n #(2, 0, 0) FANOUT_25 (c2670_wire_382, {c2670_wire_382_0, c2670_wire_382_1});
fanout_n #(2, 0, 0) FANOUT_26 (c2670_wire_386, {c2670_wire_386_0, c2670_wire_386_1});
fanout_n #(2, 0, 0) FANOUT_27 (c2670_wire_389, {c2670_wire_389_0, c2670_wire_389_1});
fanout_n #(2, 0, 0) FANOUT_28 (c2670_wire_392, {c2670_wire_392_0, c2670_wire_392_1});
fanout_n #(2, 0, 0) FANOUT_29 (c2670_wire_396, {c2670_wire_396_0, c2670_wire_396_1});
fanout_n #(2, 0, 0) FANOUT_30 (c2670_wire_401, {c2670_wire_401_0, c2670_wire_401_1});
fanout_n #(4, 0, 0) FANOUT_31 (c2670_wire_406, {c2670_wire_406_0, c2670_wire_406_1, c2670_wire_406_2, c2670_wire_406_3});
fanout_n #(3, 0, 0) FANOUT_32 (c2670_wire_428, {c2670_wire_428_0, c2670_wire_428_1, c2670_wire_428_2});
fanout_n #(2, 0, 0) FANOUT_33 (c2670_wire_416, {c2670_wire_416_0, c2670_wire_416_1});
fanout_n #(20, 0, 0) FANOUT_34 (c2670_wire_24, {c2670_wire_24_0, c2670_wire_24_1, c2670_wire_24_2, c2670_wire_24_3, c2670_wire_24_4, c2670_wire_24_5, c2670_wire_24_6, c2670_wire_24_7, c2670_wire_24_8, c2670_wire_24_9, c2670_wire_24_10, c2670_wire_24_11, c2670_wire_24_12, c2670_wire_24_13, c2670_wire_24_14, c2670_wire_24_15, c2670_wire_24_16, c2670_wire_24_17, c2670_wire_24_18, c2670_wire_24_19});
fanout_n #(6, 0, 0) FANOUT_35 (c2670_wire_13, {c2670_wire_13_0, c2670_wire_13_1, c2670_wire_13_2, c2670_wire_13_3, c2670_wire_13_4, c2670_wire_13_5});
fanout_n #(2, 0, 0) FANOUT_36 (c2670_wire_434, {c2670_wire_434_0, c2670_wire_434_1});
fanout_n #(28, 0, 0) FANOUT_37 (c2670_wire_441, {c2670_wire_441_0, c2670_wire_441_1, c2670_wire_441_2, c2670_wire_441_3, c2670_wire_441_4, c2670_wire_441_5, c2670_wire_441_6, c2670_wire_441_7, c2670_wire_441_8, c2670_wire_441_9, c2670_wire_441_10, c2670_wire_441_11, c2670_wire_441_12, c2670_wire_441_13, c2670_wire_441_14, c2670_wire_441_15, c2670_wire_441_16, c2670_wire_441_17, c2670_wire_441_18, c2670_wire_441_19, c2670_wire_441_20, c2670_wire_441_21, c2670_wire_441_22, c2670_wire_441_23, c2670_wire_441_24, c2670_wire_441_25, c2670_wire_441_26, c2670_wire_441_27});
fanout_n #(39, 0, 0) FANOUT_38 (c2670_wire_20, {c2670_wire_20_0, c2670_wire_20_1, c2670_wire_20_2, c2670_wire_20_3, c2670_wire_20_4, c2670_wire_20_5, c2670_wire_20_6, c2670_wire_20_7, c2670_wire_20_8, c2670_wire_20_9, c2670_wire_20_10, c2670_wire_20_11, c2670_wire_20_12, c2670_wire_20_13, c2670_wire_20_14, c2670_wire_20_15, c2670_wire_20_16, c2670_wire_20_17, c2670_wire_20_18, c2670_wire_20_19, c2670_wire_20_20, c2670_wire_20_21, c2670_wire_20_22, c2670_wire_20_23, c2670_wire_20_24, c2670_wire_20_25, c2670_wire_20_26, c2670_wire_20_27, c2670_wire_20_28, c2670_wire_20_29, c2670_wire_20_30, c2670_wire_20_31, c2670_wire_20_32, c2670_wire_20_33, c2670_wire_20_34, c2670_wire_20_35, c2670_wire_20_36, c2670_wire_20_37, c2670_wire_20_38});
fanout_n #(6, 0, 0) FANOUT_39 (c2670_wire_419, {c2670_wire_419_0, c2670_wire_419_1, c2670_wire_419_2, c2670_wire_419_3, c2670_wire_419_4, c2670_wire_419_5});
fanout_n #(4, 0, 0) FANOUT_40 (c2670_wire_450, {c2670_wire_450_0, c2670_wire_450_1, c2670_wire_450_2, c2670_wire_450_3});
fanout_n #(8, 0, 0) FANOUT_41 (c2670_wire_453, {c2670_wire_453_0, c2670_wire_453_1, c2670_wire_453_2, c2670_wire_453_3, c2670_wire_453_4, c2670_wire_453_5, c2670_wire_453_6, c2670_wire_453_7});
fanout_n #(2, 0, 0) FANOUT_42 (c2670_wire_464, {c2670_wire_464_0, c2670_wire_464_1});
fanout_n #(5, 0, 0) FANOUT_43 (c2670_wire_465, {c2670_wire_465_0, c2670_wire_465_1, c2670_wire_465_2, c2670_wire_465_3, c2670_wire_465_4});
fanout_n #(5, 0, 0) FANOUT_44 (c2670_wire_466, {c2670_wire_466_0, c2670_wire_466_1, c2670_wire_466_2, c2670_wire_466_3, c2670_wire_466_4});
fanout_n #(2, 0, 0) FANOUT_45 (c2670_wire_471, {c2670_wire_471_0, c2670_wire_471_1});
fanout_n #(6, 0, 0) FANOUT_46 (c2670_wire_371, {c2670_wire_371_0, c2670_wire_371_1, c2670_wire_371_2, c2670_wire_371_3, c2670_wire_371_4, c2670_wire_371_5});
fanout_n #(2, 0, 0) FANOUT_47 (c2670_wire_473, {c2670_wire_473_0, c2670_wire_473_1});
fanout_n #(5, 0, 0) FANOUT_48 (c2670_wire_483, {c2670_wire_483_0, c2670_wire_483_1, c2670_wire_483_2, c2670_wire_483_3, c2670_wire_483_4});
fanout_n #(2, 0, 0) FANOUT_49 (c2670_wire_484, {c2670_wire_484_0, c2670_wire_484_1});
fanout_n #(2, 0, 0) FANOUT_50 (c2670_wire_497, {c2670_wire_497_0, c2670_wire_497_1});
fanout_n #(7, 0, 0) FANOUT_51 (c2670_wire_489, {c2670_wire_489_0, c2670_wire_489_1, c2670_wire_489_2, c2670_wire_489_3, c2670_wire_489_4, c2670_wire_489_5, c2670_wire_489_6});
fanout_n #(5, 0, 0) FANOUT_52 (c2670_wire_525, {c2670_wire_525_0, c2670_wire_525_1, c2670_wire_525_2, c2670_wire_525_3, c2670_wire_525_4});
fanout_n #(24, 0, 0) FANOUT_53 (c2670_wire_526, {c2670_wire_526_0, c2670_wire_526_1, c2670_wire_526_2, c2670_wire_526_3, c2670_wire_526_4, c2670_wire_526_5, c2670_wire_526_6, c2670_wire_526_7, c2670_wire_526_8, c2670_wire_526_9, c2670_wire_526_10, c2670_wire_526_11, c2670_wire_526_12, c2670_wire_526_13, c2670_wire_526_14, c2670_wire_526_15, c2670_wire_526_16, c2670_wire_526_17, c2670_wire_526_18, c2670_wire_526_19, c2670_wire_526_20, c2670_wire_526_21, c2670_wire_526_22, c2670_wire_526_23});
fanout_n #(7, 0, 0) FANOUT_54 (c2670_wire_552, {c2670_wire_552_0, c2670_wire_552_1, c2670_wire_552_2, c2670_wire_552_3, c2670_wire_552_4, c2670_wire_552_5, c2670_wire_552_6});
fanout_n #(3, 0, 0) FANOUT_55 (c2670_wire_459, {c2670_wire_459_0, c2670_wire_459_1, c2670_wire_459_2});
fanout_n #(7, 0, 0) FANOUT_56 (c2670_wire_477, {c2670_wire_477_0, c2670_wire_477_1, c2670_wire_477_2, c2670_wire_477_3, c2670_wire_477_4, c2670_wire_477_5, c2670_wire_477_6});
fanout_n #(7, 0, 0) FANOUT_57 (c2670_wire_557, {c2670_wire_557_0, c2670_wire_557_1, c2670_wire_557_2, c2670_wire_557_3, c2670_wire_557_4, c2670_wire_557_5, c2670_wire_557_6});
fanout_n #(8, 0, 0) FANOUT_58 (c2670_wire_284, {c2670_wire_284_0, c2670_wire_284_1, c2670_wire_284_2, c2670_wire_284_3, c2670_wire_284_4, c2670_wire_284_5, c2670_wire_284_6, c2670_wire_284_7});
fanout_n #(9, 0, 0) FANOUT_59 (c2670_wire_302, {c2670_wire_302_0, c2670_wire_302_1, c2670_wire_302_2, c2670_wire_302_3, c2670_wire_302_4, c2670_wire_302_5, c2670_wire_302_6, c2670_wire_302_7, c2670_wire_302_8});
fanout_n #(5, 0, 0) FANOUT_60 (c2670_wire_8, {c2670_wire_8_0, c2670_wire_8_1, c2670_wire_8_2, c2670_wire_8_3, c2670_wire_8_4});
fanout_n #(3, 0, 0) FANOUT_61 (c2670_wire_571, {c2670_wire_571_0, c2670_wire_571_1, c2670_wire_571_2});
fanout_n #(7, 0, 0) FANOUT_62 (c2670_wire_329, {c2670_wire_329_0, c2670_wire_329_1, c2670_wire_329_2, c2670_wire_329_3, c2670_wire_329_4, c2670_wire_329_5, c2670_wire_329_6});
fanout_n #(8, 0, 0) FANOUT_63 (c2670_wire_347, {c2670_wire_347_0, c2670_wire_347_1, c2670_wire_347_2, c2670_wire_347_3, c2670_wire_347_4, c2670_wire_347_5, c2670_wire_347_6, c2670_wire_347_7});
fanout_n #(2, 0, 0) FANOUT_64 (c2670_wire_481, {c2670_wire_481_0, c2670_wire_481_1});
fanout_n #(6, 0, 0) FANOUT_65 (c2670_wire_574, {c2670_wire_574_0, c2670_wire_574_1, c2670_wire_574_2, c2670_wire_574_3, c2670_wire_574_4, c2670_wire_574_5});
fanout_n #(4, 0, 0) FANOUT_66 (c2670_wire_585, {c2670_wire_585_0, c2670_wire_585_1, c2670_wire_585_2, c2670_wire_585_3});
fanout_n #(7, 0, 0) FANOUT_67 (c2670_wire_586, {c2670_wire_586_0, c2670_wire_586_1, c2670_wire_586_2, c2670_wire_586_3, c2670_wire_586_4, c2670_wire_586_5, c2670_wire_586_6});
fanout_n #(2, 0, 0) FANOUT_68 (c2670_wire_587, {c2670_wire_587_0, c2670_wire_587_1});
fanout_n #(3, 0, 0) FANOUT_69 (c2670_wire_593, {c2670_wire_593_0, c2670_wire_593_1, c2670_wire_593_2});
fanout_n #(3, 0, 0) FANOUT_70 (c2670_wire_594, {c2670_wire_594_0, c2670_wire_594_1, c2670_wire_594_2});
fanout_n #(4, 0, 0) FANOUT_71 (c2670_wire_596, {c2670_wire_596_0, c2670_wire_596_1, c2670_wire_596_2, c2670_wire_596_3});
fanout_n #(5, 0, 0) FANOUT_72 (c2670_wire_597, {c2670_wire_597_0, c2670_wire_597_1, c2670_wire_597_2, c2670_wire_597_3, c2670_wire_597_4});
fanout_n #(8, 0, 0) FANOUT_73 (c2670_wire_216, {c2670_wire_216_0, c2670_wire_216_1, c2670_wire_216_2, c2670_wire_216_3, c2670_wire_216_4, c2670_wire_216_5, c2670_wire_216_6, c2670_wire_216_7});
fanout_n #(8, 0, 0) FANOUT_74 (c2670_wire_234, {c2670_wire_234_0, c2670_wire_234_1, c2670_wire_234_2, c2670_wire_234_3, c2670_wire_234_4, c2670_wire_234_5, c2670_wire_234_6, c2670_wire_234_7});
fanout_n #(4, 0, 0) FANOUT_75 (c2670_wire_255, {c2670_wire_255_0, c2670_wire_255_1, c2670_wire_255_2, c2670_wire_255_3});
fanout_n #(5, 0, 0) FANOUT_76 (c2670_wire_607, {c2670_wire_607_0, c2670_wire_607_1, c2670_wire_607_2, c2670_wire_607_3, c2670_wire_607_4});
fanout_n #(18, 0, 0) FANOUT_77 (c2670_wire_197, {c2670_wire_197_0, c2670_wire_197_1, c2670_wire_197_2, c2670_wire_197_3, c2670_wire_197_4, c2670_wire_197_5, c2670_wire_197_6, c2670_wire_197_7, c2670_wire_197_8, c2670_wire_197_9, c2670_wire_197_10, c2670_wire_197_11, c2670_wire_197_12, c2670_wire_197_13, c2670_wire_197_14, c2670_wire_197_15, c2670_wire_197_16, c2670_wire_197_17});
fanout_n #(36, 0, 0) FANOUT_78 (c2670_wire_195, {c2670_wire_195_0, c2670_wire_195_1, c2670_wire_195_2, c2670_wire_195_3, c2670_wire_195_4, c2670_wire_195_5, c2670_wire_195_6, c2670_wire_195_7, c2670_wire_195_8, c2670_wire_195_9, c2670_wire_195_10, c2670_wire_195_11, c2670_wire_195_12, c2670_wire_195_13, c2670_wire_195_14, c2670_wire_195_15, c2670_wire_195_16, c2670_wire_195_17, c2670_wire_195_18, c2670_wire_195_19, c2670_wire_195_20, c2670_wire_195_21, c2670_wire_195_22, c2670_wire_195_23, c2670_wire_195_24, c2670_wire_195_25, c2670_wire_195_26, c2670_wire_195_27, c2670_wire_195_28, c2670_wire_195_29, c2670_wire_195_30, c2670_wire_195_31, c2670_wire_195_32, c2670_wire_195_33, c2670_wire_195_34, c2670_wire_195_35});
fanout_n #(2, 0, 0) FANOUT_79 (c2670_wire_449, {c2670_wire_449_0, c2670_wire_449_1});
fanout_n #(2, 0, 0) FANOUT_80 (c2670_wire_614, {c2670_wire_614_0, c2670_wire_614_1});
fanout_n #(2, 0, 0) FANOUT_81 (c2670_wire_616, {c2670_wire_616_0, c2670_wire_616_1});
fanout_n #(2, 0, 0) FANOUT_82 (c2670_wire_523, {c2670_wire_523_0, c2670_wire_523_1});
fanout_n #(2, 0, 0) FANOUT_83 (c2670_wire_617, {c2670_wire_617_0, c2670_wire_617_1});
fanout_n #(2, 0, 0) FANOUT_84 (c2670_wire_622, {c2670_wire_622_0, c2670_wire_622_1});
fanout_n #(2, 0, 0) FANOUT_85 (c2670_wire_623, {c2670_wire_623_0, c2670_wire_623_1});
fanout_n #(2, 0, 0) FANOUT_86 (c2670_wire_624, {c2670_wire_624_0, c2670_wire_624_1});
fanout_n #(2, 0, 0) FANOUT_87 (c2670_wire_626, {c2670_wire_626_0, c2670_wire_626_1});
fanout_n #(2, 0, 0) FANOUT_88 (c2670_wire_629, {c2670_wire_629_0, c2670_wire_629_1});
fanout_n #(2, 0, 0) FANOUT_89 (c2670_wire_630, {c2670_wire_630_0, c2670_wire_630_1});
fanout_n #(2, 0, 0) FANOUT_90 (c2670_wire_632, {c2670_wire_632_0, c2670_wire_632_1});
fanout_n #(4, 0, 0) FANOUT_91 (c2670_wire_410, {c2670_wire_410_0, c2670_wire_410_1, c2670_wire_410_2, c2670_wire_410_3});
fanout_n #(4, 0, 0) FANOUT_92 (c2670_wire_634, {c2670_wire_634_0, c2670_wire_634_1, c2670_wire_634_2, c2670_wire_634_3});
fanout_n #(4, 0, 0) FANOUT_93 (c2670_wire_610, {c2670_wire_610_0, c2670_wire_610_1, c2670_wire_610_2, c2670_wire_610_3});
fanout_n #(2, 0, 0) FANOUT_94 (c2670_wire_505, {c2670_wire_505_0, c2670_wire_505_1});
fanout_n #(2, 0, 0) FANOUT_95 (c2670_wire_513, {c2670_wire_513_0, c2670_wire_513_1});
fanout_n #(4, 0, 0) FANOUT_96 (c2670_wire_716, {c2670_wire_716_0, c2670_wire_716_1, c2670_wire_716_2, c2670_wire_716_3});
fanout_n #(2, 0, 0) FANOUT_97 (c2670_wire_719, {c2670_wire_719_0, c2670_wire_719_1});
fanout_n #(2, 0, 0) FANOUT_98 (c2670_wire_518, {c2670_wire_518_0, c2670_wire_518_1});
fanout_n #(2, 0, 0) FANOUT_99 (c2670_wire_732, {c2670_wire_732_0, c2670_wire_732_1});
fanout_n #(2, 0, 0) FANOUT_100 (c2670_wire_742, {c2670_wire_742_0, c2670_wire_742_1});
fanout_n #(2, 0, 0) FANOUT_101 (c2670_wire_744, {c2670_wire_744_0, c2670_wire_744_1});
fanout_n #(3, 0, 0) FANOUT_102 (c2670_wire_755, {c2670_wire_755_0, c2670_wire_755_1, c2670_wire_755_2});
fanout_n #(2, 0, 0) FANOUT_103 (c2670_wire_758, {c2670_wire_758_0, c2670_wire_758_1});
fanout_n #(3, 0, 0) FANOUT_104 (c2670_wire_762, {c2670_wire_762_0, c2670_wire_762_1, c2670_wire_762_2});
fanout_n #(2, 0, 0) FANOUT_105 (c2670_wire_764, {c2670_wire_764_0, c2670_wire_764_1});
fanout_n #(2, 0, 0) FANOUT_106 (c2670_wire_769, {c2670_wire_769_0, c2670_wire_769_1});
fanout_n #(2, 0, 0) FANOUT_107 (c2670_wire_771, {c2670_wire_771_0, c2670_wire_771_1});
fanout_n #(2, 0, 0) FANOUT_108 (c2670_wire_452, {c2670_wire_452_0, c2670_wire_452_1});
fanout_n #(2, 0, 0) FANOUT_109 (c2670_wire_670, {c2670_wire_670_0, c2670_wire_670_1});
fanout_n #(4, 0, 0) FANOUT_110 (c2670_wire_693, {c2670_wire_693_0, c2670_wire_693_1, c2670_wire_693_2, c2670_wire_693_3});
fanout_n #(2, 0, 0) FANOUT_111 (c2670_wire_676, {c2670_wire_676_0, c2670_wire_676_1});
fanout_n #(4, 0, 0) FANOUT_112 (c2670_wire_779, {c2670_wire_779_0, c2670_wire_779_1, c2670_wire_779_2, c2670_wire_779_3});
fanout_n #(4, 0, 0) FANOUT_113 (c2670_wire_787, {c2670_wire_787_0, c2670_wire_787_1, c2670_wire_787_2, c2670_wire_787_3});
fanout_n #(4, 0, 0) FANOUT_114 (c2670_wire_792, {c2670_wire_792_0, c2670_wire_792_1, c2670_wire_792_2, c2670_wire_792_3});
fanout_n #(2, 0, 0) FANOUT_115 (c2670_wire_796, {c2670_wire_796_0, c2670_wire_796_1});
fanout_n #(4, 0, 0) FANOUT_116 (c2670_wire_805, {c2670_wire_805_0, c2670_wire_805_1, c2670_wire_805_2, c2670_wire_805_3});
fanout_n #(4, 0, 0) FANOUT_117 (c2670_wire_782, {c2670_wire_782_0, c2670_wire_782_1, c2670_wire_782_2, c2670_wire_782_3});
fanout_n #(3, 0, 0) FANOUT_118 (c2670_wire_759, {c2670_wire_759_0, c2670_wire_759_1, c2670_wire_759_2});
fanout_n #(3, 0, 0) FANOUT_119 (c2670_wire_765, {c2670_wire_765_0, c2670_wire_765_1, c2670_wire_765_2});
fanout_n #(2, 0, 0) FANOUT_120 (c2670_wire_806, {c2670_wire_806_0, c2670_wire_806_1});
fanout_n #(18, 0, 0) FANOUT_121 (c2670_wire_488, {c2670_wire_488_0, c2670_wire_488_1, c2670_wire_488_2, c2670_wire_488_3, c2670_wire_488_4, c2670_wire_488_5, c2670_wire_488_6, c2670_wire_488_7, c2670_wire_488_8, c2670_wire_488_9, c2670_wire_488_10, c2670_wire_488_11, c2670_wire_488_12, c2670_wire_488_13, c2670_wire_488_14, c2670_wire_488_15, c2670_wire_488_16, c2670_wire_488_17});
fanout_n #(2, 0, 0) FANOUT_122 (c2670_wire_827, {c2670_wire_827_0, c2670_wire_827_1});
fanout_n #(4, 0, 0) FANOUT_123 (c2670_wire_846, {c2670_wire_846_0, c2670_wire_846_1, c2670_wire_846_2, c2670_wire_846_3});
fanout_n #(2, 0, 0) FANOUT_124 (c2670_wire_850, {c2670_wire_850_0, c2670_wire_850_1});
fanout_n #(2, 0, 0) FANOUT_125 (c2670_wire_664, {c2670_wire_664_0, c2670_wire_664_1});
fanout_n #(2, 0, 0) FANOUT_126 (c2670_wire_854, {c2670_wire_854_0, c2670_wire_854_1});
fanout_n #(2, 0, 0) FANOUT_127 (c2670_wire_858, {c2670_wire_858_0, c2670_wire_858_1});
fanout_n #(2, 0, 0) FANOUT_128 (c2670_wire_862, {c2670_wire_862_0, c2670_wire_862_1});
fanout_n #(2, 0, 0) FANOUT_129 (c2670_wire_879, {c2670_wire_879_0, c2670_wire_879_1});
fanout_n #(2, 0, 0) FANOUT_130 (c2670_wire_864, {c2670_wire_864_0, c2670_wire_864_1});
fanout_n #(2, 0, 0) FANOUT_131 (c2670_wire_577, {c2670_wire_577_0, c2670_wire_577_1});
fanout_n #(3, 0, 0) FANOUT_132 (c2670_wire_899, {c2670_wire_899_0, c2670_wire_899_1, c2670_wire_899_2});
fanout_n #(2, 0, 0) FANOUT_133 (c2670_wire_928, {c2670_wire_928_0, c2670_wire_928_1});
fanout_n #(2, 0, 0) FANOUT_134 (c2670_wire_929, {c2670_wire_929_0, c2670_wire_929_1});
fanout_n #(3, 0, 0) FANOUT_135 (c2670_wire_934, {c2670_wire_934_0, c2670_wire_934_1, c2670_wire_934_2});
fanout_n #(2, 0, 0) FANOUT_136 (c2670_wire_954, {c2670_wire_954_0, c2670_wire_954_1});
fanout_n #(2, 0, 0) FANOUT_137 (c2670_wire_961, {c2670_wire_961_0, c2670_wire_961_1});
fanout_n #(2, 0, 0) FANOUT_138 (c2670_wire_963, {c2670_wire_963_0, c2670_wire_963_1});
fanout_n #(2, 0, 0) FANOUT_139 (c2670_wire_964, {c2670_wire_964_0, c2670_wire_964_1});
fanout_n #(2, 0, 0) FANOUT_140 (c2670_wire_970, {c2670_wire_970_0, c2670_wire_970_1});
fanout_n #(2, 0, 0) FANOUT_141 (c2670_wire_602, {c2670_wire_602_0, c2670_wire_602_1});
fanout_n #(2, 0, 0) FANOUT_142 (c2670_wire_604, {c2670_wire_604_0, c2670_wire_604_1});
fanout_n #(2, 0, 0) FANOUT_143 (c2670_wire_835, {c2670_wire_835_0, c2670_wire_835_1});
fanout_n #(2, 0, 0) FANOUT_144 (c2670_wire_187, {c2670_wire_187_0, c2670_wire_187_1});
fanout_n #(2, 0, 0) FANOUT_145 (c2670_wire_319, {c2670_wire_319_0, c2670_wire_319_1});
fanout_n #(2, 0, 0) FANOUT_146 (c2670_wire_955, {c2670_wire_955_0, c2670_wire_955_1});
fanout_n #(2, 0, 0) FANOUT_147 (c2670_wire_510, {c2670_wire_510_0, c2670_wire_510_1});
fanout_n #(2, 0, 0) FANOUT_148 (c2670_wire_943, {c2670_wire_943_0, c2670_wire_943_1});
fanout_n #(2, 0, 0) FANOUT_149 (c2670_wire_500, {c2670_wire_500_0, c2670_wire_500_1});
fanout_n #(2, 0, 0) FANOUT_150 (c2670_wire_939, {c2670_wire_939_0, c2670_wire_939_1});
fanout_n #(2, 0, 0) FANOUT_151 (c2670_wire_320, {c2670_wire_320_0, c2670_wire_320_1});
fanout_n #(2, 0, 0) FANOUT_152 (c2670_wire_582, {c2670_wire_582_0, c2670_wire_582_1});
fanout_n #(2, 0, 0) FANOUT_153 (c2670_wire_579, {c2670_wire_579_0, c2670_wire_579_1});
fanout_n #(2, 0, 0) FANOUT_154 (c2670_wire_580, {c2670_wire_580_0, c2670_wire_580_1});
fanout_n #(3, 0, 0) FANOUT_155 (c2670_wire_438, {c2670_wire_438_0, c2670_wire_438_1, c2670_wire_438_2});
fanout_n #(2, 0, 0) FANOUT_156 (c2670_wire_321, {c2670_wire_321_0, c2670_wire_321_1});
fanout_n #(4, 0, 0) FANOUT_157 (c2670_wire_619, {c2670_wire_619_0, c2670_wire_619_1, c2670_wire_619_2, c2670_wire_619_3});
fanout_n #(8, 0, 0) FANOUT_158 (c2670_wire_757, {c2670_wire_757_0, c2670_wire_757_1, c2670_wire_757_2, c2670_wire_757_3, c2670_wire_757_4, c2670_wire_757_5, c2670_wire_757_6, c2670_wire_757_7});
fanout_n #(2, 0, 0) FANOUT_159 (c2670_wire_945, {c2670_wire_945_0, c2670_wire_945_1});
fanout_n #(2, 0, 0) FANOUT_160 (c2670_wire_941, {c2670_wire_941_0, c2670_wire_941_1});
fanout_n #(4, 0, 0) FANOUT_161 (c2670_wire_420, {c2670_wire_420_0, c2670_wire_420_1, c2670_wire_420_2, c2670_wire_420_3});


bufg #(0, 0) BUF_1 (c2670_wire_1, G1_net_0);
bufg #(0, 0) BUF_2 (c2670_wire_2, G10_net_0);
bufg #(0, 0) BUF_3 (c2670_wire_3, G100_net_0);
or_n #(2, 0, 0) OR_1 (c2670_wire_4, {c2670_wire_5_0, c2670_wire_6});
and_n #(2, 0, 0) AND_1 (c2670_wire_7, {c2670_wire_5_1, c2670_wire_8_0});
or_n #(2, 0, 0) OR_2 (c2670_wire_5, {c2670_wire_9, c2670_wire_10});
notg #(0, 0) NOT_1 (c2670_wire_11, c2670_wire_5_2);
and_n #(2, 0, 0) AND_2 (c2670_wire_12, {c2670_wire_5_3, c2670_wire_13_0});
notg #(0, 0) NOT_2 (c2670_wire_14, c2670_wire_5_4);
and_n #(2, 0, 0) AND_3 (c2670_wire_15, {c2670_wire_5_5, c2670_wire_16});
and_n #(2, 0, 0) AND_4 (c2670_wire_17, {c2670_wire_5_6, c2670_wire_18});
and_n #(2, 0, 0) AND_5 (c2670_wire_19, {c2670_wire_20_0, c2670_wire_21});
or_n #(2, 0, 0) OR_3 (c2670_wire_22, {c2670_wire_19, c2670_wire_23});
and_n #(2, 0, 0) AND_6 (c2670_wire_9, {c2670_wire_22, c2670_wire_24_0});
and_n #(2, 0, 0) AND_7 (c2670_wire_10, {c2670_wire_25, c2670_wire_26});
notg #(0, 0) NOT_3 (c2670_wire_27, c2670_wire_20_1);
and_n #(2, 0, 0) AND_8 (c2670_wire_23, {c2670_wire_27, c2670_wire_28});
and_n #(2, 0, 0) AND_9 (c2670_wire_29, {c2670_wire_20_2, c2670_wire_30});
or_n #(2, 0, 0) OR_4 (c2670_wire_26, {c2670_wire_29, c2670_wire_31});
notg #(0, 0) NOT_4 (c2670_wire_32, c2670_wire_20_3);
and_n #(2, 0, 0) AND_10 (c2670_wire_31, {c2670_wire_32, c2670_wire_33});
notg #(0, 0) NOT_5 (c2670_wire_25, c2670_wire_24_1);
xor_n #(2, 0, 0) XOR_1 (c2670_wire_34, {c2670_wire_35_0, c2670_wire_36_0});
or_n #(2, 0, 0) OR_5 (c2670_wire_35, {c2670_wire_37, c2670_wire_38});
notg #(0, 0) NOT_6 (c2670_wire_39, c2670_wire_35_1);
or_n #(2, 0, 0) OR_6 (c2670_wire_40, {c2670_wire_35_2, c2670_wire_41});
notg #(0, 0) NOT_7 (c2670_wire_42, c2670_wire_35_3);
notg #(0, 0) NOT_8 (c2670_wire_43, c2670_wire_35_4);
notg #(0, 0) NOT_9 (c2670_wire_44, c2670_wire_35_5);
and_n #(2, 0, 0) AND_11 (c2670_wire_45, {c2670_wire_35_6, c2670_wire_46});
and_n #(2, 0, 0) AND_12 (c2670_wire_47, {c2670_wire_35_7, c2670_wire_48});
or_n #(2, 0, 0) OR_7 (c2670_wire_49, {c2670_wire_35_8, c2670_wire_50});
and_n #(2, 0, 0) AND_13 (c2670_wire_51, {c2670_wire_20_4, c2670_wire_52});
or_n #(2, 0, 0) OR_8 (c2670_wire_53, {c2670_wire_51, c2670_wire_54});
and_n #(2, 0, 0) AND_14 (c2670_wire_37, {c2670_wire_53, c2670_wire_24_2});
and_n #(2, 0, 0) AND_15 (c2670_wire_38, {c2670_wire_55, c2670_wire_56});
notg #(0, 0) NOT_10 (c2670_wire_57, c2670_wire_20_5);
and_n #(2, 0, 0) AND_16 (c2670_wire_54, {c2670_wire_57, c2670_wire_58});
and_n #(2, 0, 0) AND_17 (c2670_wire_59, {c2670_wire_20_6, c2670_wire_60});
or_n #(2, 0, 0) OR_9 (c2670_wire_56, {c2670_wire_59, c2670_wire_61});
notg #(0, 0) NOT_11 (c2670_wire_62, c2670_wire_20_7);
and_n #(2, 0, 0) AND_18 (c2670_wire_61, {c2670_wire_62, c2670_wire_63});
notg #(0, 0) NOT_12 (c2670_wire_55, c2670_wire_24_3);
and_n #(2, 0, 0) AND_19 (c2670_wire_64, {c2670_wire_3, c2670_wire_65});
bufg #(0, 0) BUF_4 (c2670_wire_66, G101_net_0);
and_n #(2, 0, 0) AND_20 (c2670_wire_67, {c2670_wire_20_8, c2670_wire_68});
or_n #(2, 0, 0) OR_10 (c2670_wire_69, {c2670_wire_67, c2670_wire_70});
notg #(0, 0) NOT_13 (c2670_wire_71, c2670_wire_20_9);
and_n #(2, 0, 0) AND_21 (c2670_wire_70, {c2670_wire_71, c2670_wire_72});
and_n #(2, 0, 0) AND_22 (c2670_wire_73, {c2670_wire_74, c2670_wire_75});
or_n #(2, 0, 0) OR_11 (c2670_wire_36, {c2670_wire_73, c2670_wire_76});
and_n #(2, 0, 0) AND_23 (c2670_wire_77, {c2670_wire_20_10, c2670_wire_78});
or_n #(2, 0, 0) OR_12 (c2670_wire_75, {c2670_wire_77, c2670_wire_79});
notg #(0, 0) NOT_14 (c2670_wire_80, c2670_wire_20_11);
and_n #(2, 0, 0) AND_24 (c2670_wire_79, {c2670_wire_80, c2670_wire_81});
notg #(0, 0) NOT_15 (c2670_wire_74, c2670_wire_24_4);
and_n #(2, 0, 0) AND_25 (c2670_wire_76, {c2670_wire_69, c2670_wire_24_5});
and_n #(2, 0, 0) AND_26 (c2670_wire_82, {c2670_wire_20_12, c2670_wire_83});
or_n #(2, 0, 0) OR_13 (c2670_wire_84, {c2670_wire_82, c2670_wire_85});
notg #(0, 0) NOT_16 (c2670_wire_86, c2670_wire_20_13);
and_n #(2, 0, 0) AND_27 (c2670_wire_85, {c2670_wire_86, c2670_wire_87});
and_n #(2, 0, 0) AND_28 (c2670_wire_88, {c2670_wire_89, c2670_wire_90});
or_n #(2, 0, 0) OR_14 (c2670_wire_91, {c2670_wire_88, c2670_wire_92});
and_n #(2, 0, 0) AND_29 (c2670_wire_93, {c2670_wire_20_14, c2670_wire_94});
or_n #(2, 0, 0) OR_15 (c2670_wire_90, {c2670_wire_93, c2670_wire_95});
notg #(0, 0) NOT_17 (c2670_wire_96, c2670_wire_20_15);
and_n #(2, 0, 0) AND_30 (c2670_wire_95, {c2670_wire_96, c2670_wire_97});
notg #(0, 0) NOT_18 (c2670_wire_89, c2670_wire_24_6);
and_n #(2, 0, 0) AND_31 (c2670_wire_92, {c2670_wire_84, c2670_wire_24_7});
and_n #(2, 0, 0) AND_32 (c2670_wire_98, {c2670_wire_66, c2670_wire_99});
bufg #(0, 0) BUF_5 (c2670_wire_100, G102_net_0);
and_n #(2, 0, 0) AND_33 (c2670_wire_101, {c2670_wire_20_16, c2670_wire_102});
or_n #(2, 0, 0) OR_16 (c2670_wire_103, {c2670_wire_101, c2670_wire_104});
notg #(0, 0) NOT_19 (c2670_wire_105, c2670_wire_20_17);
and_n #(2, 0, 0) AND_34 (c2670_wire_104, {c2670_wire_105, c2670_wire_106});
and_n #(2, 0, 0) AND_35 (c2670_wire_107, {c2670_wire_108, c2670_wire_109});
or_n #(2, 0, 0) OR_17 (c2670_wire_110, {c2670_wire_107, c2670_wire_111});
and_n #(2, 0, 0) AND_36 (c2670_wire_112, {c2670_wire_20_18, c2670_wire_113});
or_n #(2, 0, 0) OR_18 (c2670_wire_109, {c2670_wire_112, c2670_wire_114});
notg #(0, 0) NOT_20 (c2670_wire_115, c2670_wire_20_19);
and_n #(2, 0, 0) AND_37 (c2670_wire_114, {c2670_wire_115, c2670_wire_116});
notg #(0, 0) NOT_21 (c2670_wire_108, c2670_wire_24_8);
and_n #(2, 0, 0) AND_38 (c2670_wire_111, {c2670_wire_103, c2670_wire_24_9});
and_n #(2, 0, 0) AND_39 (c2670_wire_117, {c2670_wire_20_20, c2670_wire_118});
or_n #(2, 0, 0) OR_19 (c2670_wire_119, {c2670_wire_117, c2670_wire_120});
notg #(0, 0) NOT_22 (c2670_wire_121, c2670_wire_20_21);
and_n #(2, 0, 0) AND_40 (c2670_wire_120, {c2670_wire_121, c2670_wire_122});
and_n #(2, 0, 0) AND_41 (c2670_wire_123, {c2670_wire_124, c2670_wire_125});
or_n #(2, 0, 0) OR_20 (c2670_wire_126, {c2670_wire_123, c2670_wire_127});
and_n #(2, 0, 0) AND_42 (c2670_wire_128, {c2670_wire_20_22, c2670_wire_129});
or_n #(2, 0, 0) OR_21 (c2670_wire_125, {c2670_wire_128, c2670_wire_130});
notg #(0, 0) NOT_23 (c2670_wire_131, c2670_wire_20_23);
and_n #(2, 0, 0) AND_43 (c2670_wire_130, {c2670_wire_131, c2670_wire_132});
notg #(0, 0) NOT_24 (c2670_wire_124, c2670_wire_24_10);
and_n #(2, 0, 0) AND_44 (c2670_wire_127, {c2670_wire_119, c2670_wire_24_11});
and_n #(2, 0, 0) AND_45 (c2670_wire_133, {c2670_wire_100, c2670_wire_134});
bufg #(0, 0) BUF_6 (c2670_wire_135, G103_net_0);
notg #(0, 0) NOT_25 (c2670_wire_136, c2670_wire_20_24);
or_n #(2, 0, 0) OR_22 (c2670_wire_137, {c2670_wire_136, c2670_wire_138});
notg #(0, 0) NOT_26 (c2670_wire_139, c2670_wire_20_25);
and_n #(2, 0, 0) AND_46 (c2670_wire_140, {c2670_wire_139, c2670_wire_141});
and_n #(2, 0, 0) AND_47 (c2670_wire_142, {c2670_wire_20_26, c2670_wire_143});
and_n #(2, 0, 0) AND_48 (c2670_wire_144, {c2670_wire_142, c2670_wire_145});
notg #(0, 0) NOT_27 (c2670_wire_145, c2670_wire_24_12);
and_n #(2, 0, 0) AND_49 (c2670_wire_146, {c2670_wire_137, c2670_wire_24_13});
or_n #(3, 0, 0) OR_23 (c2670_wire_147, {c2670_wire_140, c2670_wire_144, c2670_wire_146});
and_n #(2, 0, 0) AND_50 (c2670_wire_148, {c2670_wire_20_27, c2670_wire_149});
or_n #(2, 0, 0) OR_24 (c2670_wire_150, {c2670_wire_148, c2670_wire_151});
notg #(0, 0) NOT_28 (c2670_wire_152, c2670_wire_20_28);
and_n #(2, 0, 0) AND_51 (c2670_wire_151, {c2670_wire_152, c2670_wire_153});
and_n #(2, 0, 0) AND_52 (c2670_wire_154, {c2670_wire_155, c2670_wire_156});
or_n #(2, 0, 0) OR_25 (c2670_wire_157, {c2670_wire_154, c2670_wire_158});
and_n #(2, 0, 0) AND_53 (c2670_wire_159, {c2670_wire_20_29, c2670_wire_160});
or_n #(2, 0, 0) OR_26 (c2670_wire_156, {c2670_wire_159, c2670_wire_161});
notg #(0, 0) NOT_29 (c2670_wire_162, c2670_wire_20_30);
and_n #(2, 0, 0) AND_54 (c2670_wire_161, {c2670_wire_162, c2670_wire_163});
notg #(0, 0) NOT_30 (c2670_wire_155, c2670_wire_24_14);
and_n #(2, 0, 0) AND_55 (c2670_wire_158, {c2670_wire_150, c2670_wire_24_15});
and_n #(2, 0, 0) AND_56 (c2670_wire_164, {c2670_wire_20_31, c2670_wire_165});
or_n #(2, 0, 0) OR_27 (c2670_wire_166, {c2670_wire_164, c2670_wire_167});
notg #(0, 0) NOT_31 (c2670_wire_168, c2670_wire_20_32);
and_n #(2, 0, 0) AND_57 (c2670_wire_167, {c2670_wire_168, c2670_wire_169});
and_n #(2, 0, 0) AND_58 (c2670_wire_170, {c2670_wire_171, c2670_wire_172});
or_n #(2, 0, 0) OR_28 (c2670_wire_173, {c2670_wire_170, c2670_wire_174});
and_n #(2, 0, 0) AND_59 (c2670_wire_175, {c2670_wire_20_33, c2670_wire_176});
or_n #(2, 0, 0) OR_29 (c2670_wire_172, {c2670_wire_175, c2670_wire_177});
notg #(0, 0) NOT_32 (c2670_wire_178, c2670_wire_20_34);
and_n #(2, 0, 0) AND_60 (c2670_wire_177, {c2670_wire_178, c2670_wire_179});
notg #(0, 0) NOT_33 (c2670_wire_171, c2670_wire_24_16);
and_n #(2, 0, 0) AND_61 (c2670_wire_174, {c2670_wire_166, c2670_wire_24_17});
notg #(0, 0) NOT_34 (c2670_wire_180, c2670_wire_181_0);
and_n #(2, 0, 0) AND_62 (c2670_wire_182, {c2670_wire_181_1, c2670_wire_183_0});
or_n #(2, 0, 0) OR_30 (c2670_wire_181, {c2670_wire_184, c2670_wire_185});
and_n #(2, 0, 0) AND_63 (c2670_wire_186, {c2670_wire_181_2, c2670_wire_187_0});
notg #(0, 0) NOT_35 (c2670_wire_188, c2670_wire_181_3);
and_n #(2, 0, 0) AND_64 (c2670_wire_189, {c2670_wire_181_4, c2670_wire_190});
and_n #(2, 0, 0) AND_65 (c2670_wire_191, {c2670_wire_181_5, c2670_wire_192});
and_n #(2, 0, 0) AND_66 (c2670_wire_193, {c2670_wire_194, c2670_wire_195_0});
or_n #(2, 0, 0) OR_31 (c2670_wire_196, {c2670_wire_193, c2670_wire_64});
and_n #(2, 0, 0) AND_67 (c2670_wire_184, {c2670_wire_196, c2670_wire_197_0});
and_n #(2, 0, 0) AND_68 (c2670_wire_185, {c2670_wire_198, c2670_wire_199});
notg #(0, 0) NOT_36 (c2670_wire_65, c2670_wire_195_1);
and_n #(2, 0, 0) AND_69 (c2670_wire_200, {c2670_wire_195_2, c2670_wire_201});
or_n #(2, 0, 0) OR_32 (c2670_wire_199, {c2670_wire_200, c2670_wire_202});
notg #(0, 0) NOT_37 (c2670_wire_203, c2670_wire_195_3);
and_n #(2, 0, 0) AND_70 (c2670_wire_202, {c2670_wire_203, c2670_wire_204});
notg #(0, 0) NOT_38 (c2670_wire_198, c2670_wire_197_1);
and_n #(2, 0, 0) AND_71 (c2670_wire_205, {c2670_wire_135, c2670_wire_206});
bufg #(0, 0) BUF_7 (c2670_wire_207, G104_net_0);
notg #(0, 0) NOT_39 (c2670_wire_208, c2670_wire_209_0);
and_n #(2, 0, 0) AND_72 (c2670_wire_210, {c2670_wire_209_1, c2670_wire_211_0});
or_n #(2, 0, 0) OR_33 (c2670_wire_209, {c2670_wire_212, c2670_wire_213});
notg #(0, 0) NOT_40 (c2670_wire_214, c2670_wire_209_2);
and_n #(2, 0, 0) AND_73 (c2670_wire_215, {c2670_wire_209_3, c2670_wire_216_0});
and_n #(2, 0, 0) AND_74 (c2670_wire_217, {c2670_wire_218, c2670_wire_195_4});
or_n #(2, 0, 0) OR_34 (c2670_wire_219, {c2670_wire_217, c2670_wire_220});
and_n #(2, 0, 0) AND_75 (c2670_wire_212, {c2670_wire_219, c2670_wire_197_2});
and_n #(2, 0, 0) AND_76 (c2670_wire_213, {c2670_wire_221, c2670_wire_222});
notg #(0, 0) NOT_41 (c2670_wire_223, c2670_wire_195_5);
and_n #(2, 0, 0) AND_77 (c2670_wire_220, {c2670_wire_223, c2670_wire_224});
and_n #(2, 0, 0) AND_78 (c2670_wire_225, {c2670_wire_195_6, c2670_wire_226});
or_n #(2, 0, 0) OR_35 (c2670_wire_222, {c2670_wire_225, c2670_wire_227});
notg #(0, 0) NOT_42 (c2670_wire_228, c2670_wire_195_7);
and_n #(2, 0, 0) AND_79 (c2670_wire_227, {c2670_wire_228, c2670_wire_229});
notg #(0, 0) NOT_43 (c2670_wire_221, c2670_wire_197_3);
notg #(0, 0) NOT_44 (c2670_wire_230, c2670_wire_211_1);
or_n #(2, 0, 0) OR_36 (c2670_wire_211, {c2670_wire_231, c2670_wire_232});
and_n #(2, 0, 0) AND_80 (c2670_wire_233, {c2670_wire_211_2, c2670_wire_234_0});
and_n #(2, 0, 0) AND_81 (c2670_wire_235, {c2670_wire_236, c2670_wire_195_8});
or_n #(2, 0, 0) OR_37 (c2670_wire_237, {c2670_wire_235, c2670_wire_238});
and_n #(2, 0, 0) AND_82 (c2670_wire_231, {c2670_wire_237, c2670_wire_197_4});
and_n #(2, 0, 0) AND_83 (c2670_wire_232, {c2670_wire_239, c2670_wire_240});
notg #(0, 0) NOT_45 (c2670_wire_241, c2670_wire_195_9);
and_n #(2, 0, 0) AND_84 (c2670_wire_238, {c2670_wire_241, c2670_wire_242});
and_n #(2, 0, 0) AND_85 (c2670_wire_243, {c2670_wire_195_10, c2670_wire_244});
or_n #(2, 0, 0) OR_38 (c2670_wire_240, {c2670_wire_243, c2670_wire_245});
notg #(0, 0) NOT_46 (c2670_wire_246, c2670_wire_195_11);
and_n #(2, 0, 0) AND_86 (c2670_wire_245, {c2670_wire_246, c2670_wire_247});
notg #(0, 0) NOT_47 (c2670_wire_239, c2670_wire_197_5);
and_n #(2, 0, 0) AND_87 (c2670_wire_248, {c2670_wire_207, c2670_wire_249});
bufg #(0, 0) BUF_8 (c2670_wire_250, G105_net_0);
or_n #(2, 0, 0) OR_39 (c2670_wire_251, {c2670_wire_252, c2670_wire_253});
and_n #(2, 0, 0) AND_88 (c2670_wire_254, {c2670_wire_251_0, c2670_wire_255_0});
and_n #(3, 0, 0) AND_89 (c2670_wire_256, {c2670_wire_251_1, c2670_wire_257, c2670_wire_258});
and_n #(2, 0, 0) AND_90 (c2670_wire_259, {c2670_wire_251_2, c2670_wire_260});
and_n #(2, 0, 0) AND_91 (c2670_wire_261, {c2670_wire_262, c2670_wire_195_12});
or_n #(2, 0, 0) OR_40 (c2670_wire_263, {c2670_wire_261, c2670_wire_264});
and_n #(2, 0, 0) AND_92 (c2670_wire_252, {c2670_wire_263, c2670_wire_197_6});
and_n #(2, 0, 0) AND_93 (c2670_wire_253, {c2670_wire_265, c2670_wire_266});
notg #(0, 0) NOT_48 (c2670_wire_267, c2670_wire_195_13);
and_n #(2, 0, 0) AND_94 (c2670_wire_264, {c2670_wire_267, c2670_wire_268});
and_n #(2, 0, 0) AND_95 (c2670_wire_269, {c2670_wire_195_14, c2670_wire_270});
or_n #(2, 0, 0) OR_41 (c2670_wire_266, {c2670_wire_269, c2670_wire_271});
notg #(0, 0) NOT_49 (c2670_wire_272, c2670_wire_195_15);
and_n #(2, 0, 0) AND_96 (c2670_wire_271, {c2670_wire_272, c2670_wire_273});
notg #(0, 0) NOT_50 (c2670_wire_265, c2670_wire_197_7);
and_n #(2, 0, 0) AND_97 (c2670_wire_274, {c2670_wire_250, c2670_wire_195_16});
bufg #(0, 0) BUF_9 (c2670_wire_275, G106_net_0);
xor_n #(2, 0, 0) XOR_2 (c2670_wire_276, {c2670_wire_277_0, c2670_wire_278});
or_n #(2, 0, 0) OR_42 (c2670_wire_277, {c2670_wire_279, c2670_wire_280});
and_n #(2, 0, 0) AND_98 (c2670_wire_281, {c2670_wire_277_1, c2670_wire_282});
and_n #(2, 0, 0) AND_99 (c2670_wire_283, {c2670_wire_277_2, c2670_wire_284_0});
or_n #(2, 0, 0) OR_43 (c2670_wire_285, {c2670_wire_274, c2670_wire_286});
and_n #(2, 0, 0) AND_100 (c2670_wire_279, {c2670_wire_285, c2670_wire_197_8});
and_n #(2, 0, 0) AND_101 (c2670_wire_280, {c2670_wire_287, c2670_wire_288});
notg #(0, 0) NOT_51 (c2670_wire_289, c2670_wire_195_17);
and_n #(2, 0, 0) AND_102 (c2670_wire_286, {c2670_wire_289, c2670_wire_290});
and_n #(2, 0, 0) AND_103 (c2670_wire_291, {c2670_wire_195_18, c2670_wire_292});
or_n #(2, 0, 0) OR_44 (c2670_wire_288, {c2670_wire_291, c2670_wire_293});
notg #(0, 0) NOT_52 (c2670_wire_294, c2670_wire_195_19);
and_n #(2, 0, 0) AND_104 (c2670_wire_293, {c2670_wire_294, c2670_wire_295});
notg #(0, 0) NOT_53 (c2670_wire_287, c2670_wire_197_9);
and_n #(2, 0, 0) AND_105 (c2670_wire_296, {c2670_wire_297_0, c2670_wire_298_0});
or_n #(2, 0, 0) OR_45 (c2670_wire_297, {c2670_wire_299, c2670_wire_300});
and_n #(2, 0, 0) AND_106 (c2670_wire_301, {c2670_wire_297_1, c2670_wire_302_0});
and_n #(2, 0, 0) AND_107 (c2670_wire_303, {c2670_wire_297_2, c2670_wire_304});
and_n #(2, 0, 0) AND_108 (c2670_wire_305, {c2670_wire_297_3, c2670_wire_306});
and_n #(2, 0, 0) AND_109 (c2670_wire_307, {c2670_wire_308, c2670_wire_195_20});
or_n #(2, 0, 0) OR_46 (c2670_wire_309, {c2670_wire_307, c2670_wire_205});
and_n #(2, 0, 0) AND_110 (c2670_wire_299, {c2670_wire_309, c2670_wire_197_10});
and_n #(2, 0, 0) AND_111 (c2670_wire_300, {c2670_wire_310, c2670_wire_311});
notg #(0, 0) NOT_54 (c2670_wire_206, c2670_wire_195_21);
and_n #(2, 0, 0) AND_112 (c2670_wire_312, {c2670_wire_195_22, c2670_wire_313});
or_n #(2, 0, 0) OR_47 (c2670_wire_311, {c2670_wire_312, c2670_wire_314});
notg #(0, 0) NOT_55 (c2670_wire_315, c2670_wire_195_23);
and_n #(2, 0, 0) AND_113 (c2670_wire_314, {c2670_wire_315, c2670_wire_316});
notg #(0, 0) NOT_56 (c2670_wire_310, c2670_wire_197_11);
notg #(0, 0) NOT_57 (c2670_wire_317, c2670_wire_275_0);
and_n #(4, 0, 0) AND_114 (c2670_wire_318, {c2670_wire_275_1, c2670_wire_319_0, c2670_wire_320_0, c2670_wire_321_0});
bufg #(0, 0) BUF_10 (c2670_wire_262, G107_net_0);
or_n #(2, 0, 0) OR_48 (c2670_wire_298, {c2670_wire_322, c2670_wire_323});
and_n #(2, 0, 0) AND_115 (c2670_wire_324, {c2670_wire_298_1, c2670_wire_325});
and_n #(2, 0, 0) AND_116 (c2670_wire_326, {c2670_wire_298_2, c2670_wire_327});
xor_n #(2, 0, 0) XOR_3 (c2670_wire_328, {c2670_wire_298_3, c2670_wire_329_0});
and_n #(2, 0, 0) AND_117 (c2670_wire_330, {c2670_wire_298_4, c2670_wire_331});
and_n #(2, 0, 0) AND_118 (c2670_wire_332, {c2670_wire_298_5, c2670_wire_333});
and_n #(2, 0, 0) AND_119 (c2670_wire_334, {c2670_wire_335, c2670_wire_195_24});
or_n #(2, 0, 0) OR_49 (c2670_wire_336, {c2670_wire_334, c2670_wire_133});
and_n #(2, 0, 0) AND_120 (c2670_wire_322, {c2670_wire_336, c2670_wire_197_12});
and_n #(2, 0, 0) AND_121 (c2670_wire_323, {c2670_wire_337, c2670_wire_338});
notg #(0, 0) NOT_58 (c2670_wire_134, c2670_wire_195_25);
and_n #(2, 0, 0) AND_122 (c2670_wire_339, {c2670_wire_195_26, c2670_wire_340});
or_n #(2, 0, 0) OR_50 (c2670_wire_338, {c2670_wire_339, c2670_wire_341});
notg #(0, 0) NOT_59 (c2670_wire_342, c2670_wire_195_27);
and_n #(2, 0, 0) AND_123 (c2670_wire_341, {c2670_wire_342, c2670_wire_343});
notg #(0, 0) NOT_60 (c2670_wire_337, c2670_wire_197_13);
or_n #(2, 0, 0) OR_51 (c2670_wire_183, {c2670_wire_344, c2670_wire_345});
and_n #(2, 0, 0) AND_124 (c2670_wire_346, {c2670_wire_183_1, c2670_wire_347_0});
and_n #(2, 0, 0) AND_125 (c2670_wire_348, {c2670_wire_349, c2670_wire_195_28});
or_n #(2, 0, 0) OR_52 (c2670_wire_350, {c2670_wire_348, c2670_wire_98});
and_n #(2, 0, 0) AND_126 (c2670_wire_344, {c2670_wire_350, c2670_wire_197_14});
and_n #(2, 0, 0) AND_127 (c2670_wire_345, {c2670_wire_351, c2670_wire_352});
notg #(0, 0) NOT_61 (c2670_wire_99, c2670_wire_195_29);
and_n #(2, 0, 0) AND_128 (c2670_wire_353, {c2670_wire_195_30, c2670_wire_354});
or_n #(2, 0, 0) OR_53 (c2670_wire_352, {c2670_wire_353, c2670_wire_355});
notg #(0, 0) NOT_62 (c2670_wire_356, c2670_wire_195_31);
and_n #(2, 0, 0) AND_129 (c2670_wire_355, {c2670_wire_356, c2670_wire_357});
notg #(0, 0) NOT_63 (c2670_wire_351, c2670_wire_197_15);
or_n #(2, 0, 0) OR_54 (c2670_wire_278, {c2670_wire_358, c2670_wire_359});
and_n #(2, 0, 0) AND_130 (c2670_wire_360, {c2670_wire_361, c2670_wire_195_32});
or_n #(2, 0, 0) OR_55 (c2670_wire_362, {c2670_wire_360, c2670_wire_248});
and_n #(2, 0, 0) AND_131 (c2670_wire_358, {c2670_wire_362, c2670_wire_197_16});
and_n #(2, 0, 0) AND_132 (c2670_wire_359, {c2670_wire_363, c2670_wire_364});
notg #(0, 0) NOT_64 (c2670_wire_249, c2670_wire_195_33);
and_n #(2, 0, 0) AND_133 (c2670_wire_365, {c2670_wire_195_34, c2670_wire_366});
or_n #(2, 0, 0) OR_56 (c2670_wire_364, {c2670_wire_365, c2670_wire_367});
notg #(0, 0) NOT_65 (c2670_wire_368, c2670_wire_195_35);
and_n #(2, 0, 0) AND_134 (c2670_wire_367, {c2670_wire_368, c2670_wire_369});
notg #(0, 0) NOT_66 (c2670_wire_363, c2670_wire_197_17);
bufg #(0, 0) BUF_11 (c2670_wire_236, G108_net_0);
xor_n #(2, 0, 0) XOR_4 (c2670_wire_370, {c2670_wire_371_0, c2670_wire_372});
and_n #(2, 0, 0) AND_135 (c2670_wire_373, {c2670_wire_370_0, c2670_wire_374});
or_n #(2, 0, 0) OR_57 (c2670_wire_375, {c2670_wire_376, c2670_wire_377});
xor_n #(2, 0, 0) XOR_5 (c2670_wire_374, {c2670_wire_375_0, c2670_wire_378_0});
xor_n #(2, 0, 0) XOR_6 (c2670_wire_379, {c2670_wire_375_1, c2670_wire_378_1});
bufg #(0, 0) BUF_12 (c2670_wire_218, G109_net_0);
or_n #(2, 0, 0) OR_58 (c2670_wire_378, {c2670_wire_380, c2670_wire_381});
xor_n #(2, 0, 0) XOR_7 (c2670_wire_382, {c2670_wire_329_1, c2670_wire_383});
and_n #(2, 0, 0) AND_136 (c2670_wire_384, {c2670_wire_382_0, c2670_wire_385});
and_n #(2, 0, 0) AND_137 (c2670_wire_386, {c2670_wire_2, c2670_wire_387});
bufg #(0, 0) BUF_13 (c2670_wire_388, G11_net_0);
bufg #(0, 0) BUF_14 (c2670_wire_194, G110_net_0);
or_n #(2, 0, 0) OR_59 (c2670_wire_389, {c2670_wire_390, c2670_wire_391});
xor_n #(2, 0, 0) XOR_8 (c2670_wire_385, {c2670_wire_389_0, c2670_wire_392_0});
xor_n #(2, 0, 0) XOR_9 (c2670_wire_393, {c2670_wire_389_1, c2670_wire_392_1});
or_n #(2, 0, 0) OR_60 (c2670_wire_392, {c2670_wire_394, c2670_wire_395});
bufg #(0, 0) BUF_15 (c2670_wire_349, G111_net_0);
or_n #(2, 0, 0) OR_61 (c2670_wire_396, {c2670_wire_397, c2670_wire_398});
and_n #(2, 0, 0) AND_138 (c2670_wire_399, {c2670_wire_396_0, c2670_wire_400});
or_n #(2, 0, 0) OR_62 (c2670_wire_401, {c2670_wire_402, c2670_wire_403});
and_n #(2, 0, 0) AND_139 (c2670_wire_404, {c2670_wire_401_0, c2670_wire_405});
or_n #(2, 0, 0) OR_63 (c2670_wire_406, {c2670_wire_407, c2670_wire_408});
and_n #(2, 0, 0) AND_140 (c2670_wire_409, {c2670_wire_406_0, c2670_wire_410_0});
and_n #(2, 0, 0) AND_141 (c2670_wire_411, {c2670_wire_406_1, c2670_wire_410_1});
notg #(0, 0) NOT_67 (c2670_wire_412, c2670_wire_413);
and_n #(2, 0, 0) AND_142 (c2670_wire_413, {c2670_wire_414, c2670_wire_415});
and_n #(2, 0, 0) AND_143 (c2670_wire_414, {c2670_wire_416_0, c2670_wire_417});
notg #(0, 0) NOT_68 (c2670_wire_418, c2670_wire_419_0);
and_n #(2, 0, 0) AND_144 (c2670_wire_415, {c2670_wire_418, c2670_wire_420_0});
notg #(0, 0) NOT_69 (c2670_wire_421, c2670_wire_422);
and_n #(2, 0, 0) AND_145 (c2670_wire_422, {c2670_wire_423, c2670_wire_424});
and_n #(2, 0, 0) AND_146 (c2670_wire_423, {c2670_wire_416_1, c2670_wire_420_1});
nand_n #(2, 0, 0) NAND_1 (c2670_wire_425, {c2670_wire_1, c2670_wire_426});
notg #(0, 0) NOT_70 (c2670_wire_427, c2670_wire_419_1);
and_n #(2, 0, 0) AND_147 (c2670_wire_424, {c2670_wire_427, c2670_wire_425});
bufg #(0, 0) BUF_16 (c2670_wire_335, G112_net_0);
bufg #(0, 0) BUF_17 (c2670_wire_308, G113_net_0);
bufg #(0, 0) BUF_18 (c2670_wire_361, G114_net_0);
bufg #(0, 0) BUF_19 (c2670_wire_428, G115_net_0);
bufg #(0, 0) BUF_20 (c2670_wire_416, G116_net_0);
bufg #(0, 0) BUF_21 (c2670_wire_24, G117_net_0);
notg #(0, 0) NOT_71 (c2670_wire_429, c2670_wire_24_18);
and_n #(2, 0, 0) AND_148 (c2670_wire_430, {c2670_wire_24_19, c2670_wire_431});
bufg #(0, 0) BUF_22 (c2670_wire_13, G118_net_0);
notg #(0, 0) NOT_72 (c2670_wire_41, c2670_wire_13_1);
notg #(0, 0) NOT_73 (c2670_wire_432, c2670_wire_13_2);
and_n #(2, 0, 0) AND_149 (c2670_wire_50, {c2670_wire_13_3, c2670_wire_433});
bufg #(0, 0) BUF_23 (c2670_wire_434, G119_net_0);
and_n #(2, 0, 0) AND_150 (c2670_wire_435, {c2670_wire_434_0, c2670_wire_436});
and_n #(3, 0, 0) AND_151 (c2670_wire_437, {c2670_wire_434_1, c2670_wire_419_2, c2670_wire_438_0});
and_n #(3, 0, 0) AND_152 (c2670_wire_439, {c2670_wire_388, c2670_wire_419_3, c2670_wire_440});
bufg #(0, 0) BUF_24 (c2670_wire_441, G12_net_0);
bufg #(0, 0) BUF_25 (c2670_wire_20, G120_net_0);
and_n #(2, 0, 0) AND_153 (c2670_wire_442, {c2670_wire_20_35, c2670_wire_443});
notg #(0, 0) NOT_74 (c2670_wire_444, c2670_wire_20_36);
and_n #(2, 0, 0) AND_154 (c2670_wire_445, {c2670_wire_20_37, c2670_wire_446});
notg #(0, 0) NOT_75 (c2670_wire_447, c2670_wire_20_38);
bufg #(0, 0) BUF_26 (c2670_wire_419, G121_net_0);
and_n #(3, 0, 0) AND_155 (c2670_wire_448, {c2670_wire_419_4, c2670_wire_449_0, c2670_wire_438_1});
bufg #(0, 0) BUF_27 (c2670_wire_450, G122_net_0);
notg #(0, 0) NOT_76 (c2670_wire_6, c2670_wire_450_0);
or_n #(2, 0, 0) OR_64 (c2670_wire_451, {c2670_wire_450_1, c2670_wire_452_0});
notg #(0, 0) NOT_77 (c2670_wire_433, c2670_wire_450_2);
bufg #(0, 0) BUF_28 (c2670_wire_453, G123_net_0);
notg #(0, 0) NOT_78 (c2670_wire_454, c2670_wire_453_0);
and_n #(2, 0, 0) AND_156 (c2670_wire_455, {c2670_wire_453_1, c2670_wire_456});
and_n #(2, 0, 0) AND_157 (c2670_wire_457, {c2670_wire_453_2, c2670_wire_91_0});
and_n #(2, 0, 0) AND_158 (c2670_wire_458, {c2670_wire_453_3, c2670_wire_459_0});
notg #(0, 0) NOT_79 (c2670_wire_460, c2670_wire_453_4);
and_n #(2, 0, 0) AND_159 (c2670_wire_461, {c2670_wire_453_5, c2670_wire_462});
bufg #(0, 0) BUF_29 (c2670_wire_463, G124_net_0);
notg #(0, 0) NOT_80 (c2670_wire_464, c2670_wire_463);
bufg #(0, 0) BUF_30 (c2670_wire_465, G125_net_0);
and_n #(2, 0, 0) AND_160 (c2670_wire_397, {c2670_wire_465_0, c2670_wire_466_0});
and_n #(2, 0, 0) AND_161 (c2670_wire_467, {c2670_wire_465_1, c2670_wire_468});
bufg #(0, 0) BUF_31 (c2670_wire_466, G126_net_0);
and_n #(2, 0, 0) AND_162 (c2670_wire_469, {c2670_wire_466_1, c2670_wire_470});
bufg #(0, 0) BUF_32 (c2670_wire_471, G127_net_0);
or_n #(2, 0, 0) OR_65 (c2670_wire_472, {c2670_wire_471_0, c2670_wire_188});
bufg #(0, 0) BUF_33 (c2670_wire_371, G128_net_0);
or_n #(2, 0, 0) OR_66 (c2670_wire_473, {c2670_wire_474, c2670_wire_475});
and_n #(2, 0, 0) AND_163 (c2670_wire_476, {c2670_wire_473_0, c2670_wire_477_0});
and_n #(2, 0, 0) AND_164 (c2670_wire_474, {c2670_wire_441_0, c2670_wire_478});
notg #(0, 0) NOT_81 (c2670_wire_479, c2670_wire_441_1);
and_n #(2, 0, 0) AND_165 (c2670_wire_475, {c2670_wire_479, c2670_wire_157_0});
and_n #(2, 0, 0) AND_166 (c2670_wire_480, {c2670_wire_371_1, c2670_wire_481_0});
and_n #(2, 0, 0) AND_167 (c2670_wire_482, {c2670_wire_371_2, c2670_wire_36_1});
bufg #(0, 0) BUF_34 (c2670_wire_483, G129_net_0);
or_n #(2, 0, 0) OR_67 (c2670_wire_484, {c2670_wire_485, c2670_wire_281});
and_n #(2, 0, 0) AND_168 (c2670_wire_486, {c2670_wire_484_0, c2670_wire_284_1});
and_n #(2, 0, 0) AND_169 (c2670_wire_485, {c2670_wire_487, c2670_wire_488_0});
notg #(0, 0) NOT_82 (c2670_wire_282, c2670_wire_488_1);
and_n #(2, 0, 0) AND_170 (c2670_wire_376, {c2670_wire_483_0, c2670_wire_489_0});
and_n #(2, 0, 0) AND_171 (c2670_wire_490, {c2670_wire_483_1, c2670_wire_491});
notg #(0, 0) NOT_83 (c2670_wire_492, c2670_wire_441_2);
and_n #(3, 0, 0) AND_172 (c2670_wire_493, {c2670_wire_441_3, c2670_wire_494, c2670_wire_495});
and_n #(2, 0, 0) AND_173 (c2670_wire_496, {c2670_wire_441_4, c2670_wire_497_0});
notg #(0, 0) NOT_84 (c2670_wire_16, c2670_wire_441_5);
and_n #(2, 0, 0) AND_174 (c2670_wire_498, {c2670_wire_441_6, c2670_wire_497_1});
notg #(0, 0) NOT_85 (c2670_wire_18, c2670_wire_441_7);
and_n #(2, 0, 0) AND_175 (c2670_wire_499, {c2670_wire_441_8, c2670_wire_500_0});
notg #(0, 0) NOT_86 (c2670_wire_501, c2670_wire_441_9);
and_n #(2, 0, 0) AND_176 (c2670_wire_502, {c2670_wire_441_10, c2670_wire_500_1});
notg #(0, 0) NOT_87 (c2670_wire_503, c2670_wire_441_11);
and_n #(2, 0, 0) AND_177 (c2670_wire_504, {c2670_wire_441_12, c2670_wire_505_0});
notg #(0, 0) NOT_88 (c2670_wire_506, c2670_wire_441_13);
and_n #(2, 0, 0) AND_178 (c2670_wire_507, {c2670_wire_441_14, c2670_wire_505_1});
notg #(0, 0) NOT_89 (c2670_wire_508, c2670_wire_441_15);
and_n #(2, 0, 0) AND_179 (c2670_wire_509, {c2670_wire_441_16, c2670_wire_510_0});
notg #(0, 0) NOT_90 (c2670_wire_46, c2670_wire_441_17);
and_n #(2, 0, 0) AND_180 (c2670_wire_511, {c2670_wire_441_18, c2670_wire_510_1});
notg #(0, 0) NOT_91 (c2670_wire_48, c2670_wire_441_19);
and_n #(2, 0, 0) AND_181 (c2670_wire_512, {c2670_wire_441_20, c2670_wire_513_0});
notg #(0, 0) NOT_92 (c2670_wire_514, c2670_wire_441_21);
and_n #(2, 0, 0) AND_182 (c2670_wire_515, {c2670_wire_441_22, c2670_wire_513_1});
notg #(0, 0) NOT_93 (c2670_wire_516, c2670_wire_441_23);
and_n #(2, 0, 0) AND_183 (c2670_wire_517, {c2670_wire_441_24, c2670_wire_518_0});
notg #(0, 0) NOT_94 (c2670_wire_519, c2670_wire_441_25);
and_n #(2, 0, 0) AND_184 (c2670_wire_520, {c2670_wire_441_26, c2670_wire_518_1});
notg #(0, 0) NOT_95 (c2670_wire_521, c2670_wire_441_27);
bufg #(0, 0) BUF_35 (c2670_wire_497, G13_net_0);
bufg #(0, 0) BUF_36 (c2670_wire_489, G130_net_0);
and_n #(2, 0, 0) AND_185 (c2670_wire_522, {c2670_wire_489_1, c2670_wire_523_0});
and_n #(2, 0, 0) AND_186 (c2670_wire_524, {c2670_wire_489_2, c2670_wire_110_0});
bufg #(0, 0) BUF_37 (c2670_wire_525, G131_net_0);
and_n #(2, 0, 0) AND_187 (c2670_wire_526, {c2670_wire_186, c2670_wire_527});
and_n #(2, 0, 0) AND_188 (c2670_wire_528, {c2670_wire_526_0, c2670_wire_529});
and_n #(2, 0, 0) AND_189 (c2670_wire_530, {c2670_wire_526_1, c2670_wire_531});
and_n #(2, 0, 0) AND_190 (c2670_wire_532, {c2670_wire_526_2, c2670_wire_533});
and_n #(2, 0, 0) AND_191 (c2670_wire_534, {c2670_wire_526_3, c2670_wire_535});
and_n #(2, 0, 0) AND_192 (c2670_wire_536, {c2670_wire_526_4, c2670_wire_537});
and_n #(2, 0, 0) AND_193 (c2670_wire_538, {c2670_wire_526_5, c2670_wire_539});
notg #(0, 0) NOT_96 (c2670_wire_540, c2670_wire_526_6);
notg #(0, 0) NOT_97 (c2670_wire_541, c2670_wire_526_7);
notg #(0, 0) NOT_98 (c2670_wire_542, c2670_wire_526_8);
notg #(0, 0) NOT_99 (c2670_wire_543, c2670_wire_526_9);
and_n #(2, 0, 0) AND_194 (c2670_wire_544, {c2670_wire_526_10, c2670_wire_545});
and_n #(2, 0, 0) AND_195 (c2670_wire_546, {c2670_wire_526_11, c2670_wire_547});
notg #(0, 0) NOT_100 (c2670_wire_548, c2670_wire_526_12);
notg #(0, 0) NOT_101 (c2670_wire_549, c2670_wire_526_13);
notg #(0, 0) NOT_102 (c2670_wire_550, c2670_wire_526_14);
notg #(0, 0) NOT_103 (c2670_wire_551, c2670_wire_526_15);
nor_n #(2, 0, 0) NOR_1 (c2670_wire_527, {c2670_wire_209_4, c2670_wire_471_1});
and_n #(2, 0, 0) AND_196 (c2670_wire_380, {c2670_wire_525_0, c2670_wire_552_0});
and_n #(2, 0, 0) AND_197 (c2670_wire_553, {c2670_wire_525_1, c2670_wire_554});
bufg #(0, 0) BUF_38 (c2670_wire_552, G132_net_0);
nor_n #(2, 0, 0) NOR_2 (c2670_wire_459, {c2670_wire_13_4, c2670_wire_35_9});
and_n #(2, 0, 0) AND_198 (c2670_wire_555, {c2670_wire_552_1, c2670_wire_556});
bufg #(0, 0) BUF_39 (c2670_wire_477, G133_net_0);
and_n #(2, 0, 0) AND_199 (c2670_wire_407, {c2670_wire_477_1, c2670_wire_557_0});
notg #(0, 0) NOT_104 (c2670_wire_558, c2670_wire_477_2);
notg #(0, 0) NOT_105 (c2670_wire_559, c2670_wire_477_3);
bufg #(0, 0) BUF_40 (c2670_wire_557, G134_net_0);
notg #(0, 0) NOT_106 (c2670_wire_560, c2670_wire_557_1);
notg #(0, 0) NOT_107 (c2670_wire_561, c2670_wire_557_2);
xor_n #(2, 0, 0) XOR_10 (c2670_wire_562, {c2670_wire_557_3, c2670_wire_173_0});
and_n #(2, 0, 0) AND_200 (c2670_wire_563, {c2670_wire_557_4, c2670_wire_564});
bufg #(0, 0) BUF_41 (c2670_wire_284, G135_net_0);
and_n #(2, 0, 0) AND_201 (c2670_wire_402, {c2670_wire_284_2, c2670_wire_302_1});
bufg #(0, 0) BUF_42 (c2670_wire_302, G136_net_0);
notg #(0, 0) NOT_108 (c2670_wire_537, c2670_wire_302_2);
and_n #(2, 0, 0) AND_202 (c2670_wire_565, {c2670_wire_302_3, c2670_wire_566});
bufg #(0, 0) BUF_43 (c2670_wire_567, G137_net_0);
or_n #(2, 0, 0) OR_68 (c2670_wire_8, {c2670_wire_568, c2670_wire_430});
and_n #(2, 0, 0) AND_203 (c2670_wire_569, {c2670_wire_8_1, c2670_wire_451});
and_n #(2, 0, 0) AND_204 (c2670_wire_570, {c2670_wire_8_2, c2670_wire_460});
notg #(0, 0) NOT_109 (c2670_wire_571, c2670_wire_567);
bufg #(0, 0) BUF_44 (c2670_wire_329, G138_net_0);
notg #(0, 0) NOT_110 (c2670_wire_529, c2670_wire_329_2);
notg #(0, 0) NOT_111 (c2670_wire_325, c2670_wire_329_3);
notg #(0, 0) NOT_112 (c2670_wire_327, c2670_wire_329_4);
and_n #(2, 0, 0) AND_205 (c2670_wire_572, {c2670_wire_329_5, c2670_wire_573});
bufg #(0, 0) BUF_45 (c2670_wire_347, G139_net_0);
and_n #(2, 0, 0) AND_206 (c2670_wire_390, {c2670_wire_347_1, c2670_wire_574_0});
and_n #(4, 0, 0) AND_207 (c2670_wire_575, {c2670_wire_347_2, c2670_wire_574_1, c2670_wire_216_1, c2670_wire_234_1});
notg #(0, 0) NOT_113 (c2670_wire_531, c2670_wire_347_3);
and_n #(2, 0, 0) AND_208 (c2670_wire_576, {c2670_wire_347_4, c2670_wire_577_0});
bufg #(0, 0) BUF_46 (c2670_wire_481, G14_net_0);
bufg #(0, 0) BUF_47 (c2670_wire_574, G140_net_0);
xor_n #(2, 0, 0) XOR_11 (c2670_wire_578, {c2670_wire_579_0, c2670_wire_580_0});
and_n #(2, 0, 0) AND_209 (c2670_wire_581, {c2670_wire_578, c2670_wire_582_0});
nor_n #(2, 0, 0) NOR_3 (c2670_wire_583, {c2670_wire_582_1, c2670_wire_584});
xor_n #(2, 0, 0) XOR_12 (c2670_wire_584, {c2670_wire_579_1, c2670_wire_580_1});
or_n #(2, 0, 0) OR_69 (c2670_wire_585, {c2670_wire_581, c2670_wire_583});
and_n #(3, 0, 0) AND_210 (c2670_wire_586, {c2670_wire_214, c2670_wire_472, c2670_wire_187_1});
and_n #(3, 0, 0) AND_211 (c2670_wire_587, {c2670_wire_586_0, c2670_wire_540, c2670_wire_588});
and_n #(3, 0, 0) AND_212 (c2670_wire_589, {c2670_wire_586_1, c2670_wire_590, c2670_wire_542});
and_n #(2, 0, 0) AND_213 (c2670_wire_591, {c2670_wire_586_2, c2670_wire_592});
and_n #(3, 0, 0) AND_214 (c2670_wire_593, {c2670_wire_586_3, c2670_wire_562, c2670_wire_548});
and_n #(3, 0, 0) AND_215 (c2670_wire_594, {c2670_wire_586_4, c2670_wire_549, c2670_wire_595});
and_n #(3, 0, 0) AND_216 (c2670_wire_596, {c2670_wire_586_5, c2670_wire_328, c2670_wire_550});
and_n #(3, 0, 0) AND_217 (c2670_wire_597, {c2670_wire_586_6, c2670_wire_551, c2670_wire_598});
notg #(0, 0) NOT_114 (c2670_wire_533, c2670_wire_574_2);
and_n #(2, 0, 0) AND_218 (c2670_wire_599, {c2670_wire_574_3, c2670_wire_600});
bufg #(0, 0) BUF_48 (c2670_wire_216, G141_net_0);
and_n #(2, 0, 0) AND_219 (c2670_wire_394, {c2670_wire_216_2, c2670_wire_234_2});
notg #(0, 0) NOT_115 (c2670_wire_539, c2670_wire_216_3);
and_n #(2, 0, 0) AND_220 (c2670_wire_601, {c2670_wire_216_4, c2670_wire_602_0});
bufg #(0, 0) BUF_49 (c2670_wire_234, G142_net_0);
notg #(0, 0) NOT_116 (c2670_wire_535, c2670_wire_234_3);
and_n #(2, 0, 0) AND_221 (c2670_wire_603, {c2670_wire_234_4, c2670_wire_604_0});
bufg #(0, 0) BUF_50 (c2670_wire_255, G143_net_0);
and_n #(2, 0, 0) AND_222 (c2670_wire_605, {c2670_wire_255_1, c2670_wire_606});
bufg #(0, 0) BUF_51 (c2670_wire_607, G144_net_0);
or_n #(2, 0, 0) OR_70 (c2670_wire_608, {c2670_wire_607_0, c2670_wire_254});
and_n #(2, 0, 0) AND_223 (c2670_wire_609, {c2670_wire_607_1, c2670_wire_610_0});
and_n #(2, 0, 0) AND_224 (c2670_wire_611, {c2670_wire_607_2, c2670_wire_610_1});
bufg #(0, 0) BUF_52 (c2670_wire_197, G145_net_0);
bufg #(0, 0) BUF_53 (c2670_wire_195, G146_net_0);
bufg #(0, 0) BUF_54 (c2670_wire_449, G147_net_0);
notg #(0, 0) NOT_117 (c2670_wire_612, c2670_wire_459_1);
notg #(0, 0) NOT_118 (c2670_wire_613, c2670_wire_449_1);
bufg #(0, 0) BUF_55 (c2670_wire_614, G148_net_0);
and_n #(2, 0, 0) AND_225 (c2670_wire_615, {c2670_wire_614_0, c2670_wire_616_0});
bufg #(0, 0) BUF_56 (c2670_wire_616, G149_net_0);
bufg #(0, 0) BUF_57 (c2670_wire_523, G15_net_0);
bufg #(0, 0) BUF_58 (c2670_wire_617, G150_net_0);
and_n #(2, 0, 0) AND_226 (c2670_wire_618, {c2670_wire_585_0, c2670_wire_619_0});
and_n #(2, 0, 0) AND_227 (c2670_wire_620, {c2670_wire_585_1, c2670_wire_619_1});
and_n #(2, 0, 0) AND_228 (c2670_wire_621, {c2670_wire_617_0, c2670_wire_622_0});
bufg #(0, 0) BUF_59 (c2670_wire_622, G151_net_0);
bufg #(0, 0) BUF_60 (c2670_wire_623, G152_net_0);
or_n #(2, 0, 0) OR_71 (c2670_wire_624, {c2670_wire_296, c2670_wire_625});
nor_n #(2, 0, 0) NOR_4 (c2670_wire_625, {c2670_wire_297_4, c2670_wire_298_6});
or_n #(2, 0, 0) OR_72 (c2670_wire_626, {c2670_wire_182, c2670_wire_627});
nor_n #(2, 0, 0) NOR_5 (c2670_wire_627, {c2670_wire_183_2, c2670_wire_181_6});
and_n #(2, 0, 0) AND_229 (c2670_wire_628, {c2670_wire_623_0, c2670_wire_629_0});
bufg #(0, 0) BUF_61 (c2670_wire_629, G153_net_0);
bufg #(0, 0) BUF_62 (c2670_wire_630, G154_net_0);
and_n #(2, 0, 0) AND_230 (c2670_wire_631, {c2670_wire_630_0, c2670_wire_632_0});
bufg #(0, 0) BUF_63 (c2670_wire_632, G155_net_0);
bufg #(0, 0) BUF_64 (c2670_wire_372, G156_net_0);
bufg #(0, 0) BUF_65 (c2670_wire_383, G157_net_0);
nor_n #(2, 0, 0) NOR_6 (c2670_wire_633, {c2670_wire_370_1, c2670_wire_379});
or_n #(2, 0, 0) OR_73 (c2670_wire_410, {c2670_wire_373, c2670_wire_633});
or_n #(2, 0, 0) OR_74 (c2670_wire_634, {c2670_wire_210, c2670_wire_635});
nor_n #(2, 0, 0) NOR_7 (c2670_wire_635, {c2670_wire_209_5, c2670_wire_211_3});
nor_n #(2, 0, 0) NOR_8 (c2670_wire_636, {c2670_wire_382_1, c2670_wire_393});
or_n #(2, 0, 0) OR_75 (c2670_wire_610, {c2670_wire_384, c2670_wire_636});
bufg #(0, 0) BUF_66 (c2670_wire_505, G16_net_0);
or_n #(2, 0, 0) OR_76 (c2670_wire_468, {c2670_wire_496, c2670_wire_15});
nor_n #(2, 0, 0) NOR_9 (c2670_wire_637, {c2670_wire_638, c2670_wire_465_2});
or_n #(2, 0, 0) OR_77 (c2670_wire_639, {c2670_wire_637, c2670_wire_467});
or_n #(2, 0, 0) OR_78 (c2670_wire_638, {c2670_wire_498, c2670_wire_17});
or_n #(2, 0, 0) OR_79 (c2670_wire_470, {c2670_wire_509, c2670_wire_45});
nor_n #(2, 0, 0) NOR_10 (c2670_wire_640, {c2670_wire_641, c2670_wire_466_2});
or_n #(2, 0, 0) OR_80 (c2670_wire_642, {c2670_wire_640, c2670_wire_469});
or_n #(2, 0, 0) OR_81 (c2670_wire_641, {c2670_wire_511, c2670_wire_47});
or_n #(2, 0, 0) OR_82 (c2670_wire_491, {c2670_wire_499, c2670_wire_643});
and_n #(2, 0, 0) AND_231 (c2670_wire_643, {c2670_wire_501, c2670_wire_91_1});
nor_n #(2, 0, 0) NOR_11 (c2670_wire_644, {c2670_wire_645, c2670_wire_483_2});
or_n #(2, 0, 0) OR_83 (c2670_wire_646, {c2670_wire_644, c2670_wire_490});
or_n #(2, 0, 0) OR_84 (c2670_wire_645, {c2670_wire_502, c2670_wire_647});
and_n #(2, 0, 0) AND_232 (c2670_wire_647, {c2670_wire_503, c2670_wire_91_2});
or_n #(2, 0, 0) OR_85 (c2670_wire_554, {c2670_wire_504, c2670_wire_648});
and_n #(2, 0, 0) AND_233 (c2670_wire_648, {c2670_wire_506, c2670_wire_126_0});
nor_n #(2, 0, 0) NOR_12 (c2670_wire_649, {c2670_wire_650, c2670_wire_525_2});
or_n #(2, 0, 0) OR_86 (c2670_wire_651, {c2670_wire_649, c2670_wire_553});
or_n #(2, 0, 0) OR_87 (c2670_wire_650, {c2670_wire_507, c2670_wire_652});
and_n #(2, 0, 0) AND_234 (c2670_wire_652, {c2670_wire_508, c2670_wire_126_1});
or_n #(2, 0, 0) OR_88 (c2670_wire_556, {c2670_wire_512, c2670_wire_653});
and_n #(2, 0, 0) AND_235 (c2670_wire_653, {c2670_wire_514, c2670_wire_147_0});
nor_n #(2, 0, 0) NOR_13 (c2670_wire_654, {c2670_wire_655, c2670_wire_552_2});
or_n #(2, 0, 0) OR_89 (c2670_wire_656, {c2670_wire_654, c2670_wire_555});
or_n #(2, 0, 0) OR_90 (c2670_wire_655, {c2670_wire_515, c2670_wire_657});
and_n #(2, 0, 0) AND_236 (c2670_wire_657, {c2670_wire_516, c2670_wire_147_1});
or_n #(2, 0, 0) OR_91 (c2670_wire_564, {c2670_wire_517, c2670_wire_658});
and_n #(2, 0, 0) AND_237 (c2670_wire_658, {c2670_wire_519, c2670_wire_173_1});
nor_n #(2, 0, 0) NOR_14 (c2670_wire_659, {c2670_wire_660, c2670_wire_557_5});
or_n #(2, 0, 0) OR_92 (c2670_wire_661, {c2670_wire_659, c2670_wire_563});
or_n #(2, 0, 0) OR_93 (c2670_wire_660, {c2670_wire_520, c2670_wire_662});
and_n #(2, 0, 0) AND_238 (c2670_wire_662, {c2670_wire_521, c2670_wire_173_2});
and_n #(2, 0, 0) AND_239 (c2670_wire_663, {c2670_wire_488_2, c2670_wire_664_0});
or_n #(2, 0, 0) OR_94 (c2670_wire_566, {c2670_wire_663, c2670_wire_303});
notg #(0, 0) NOT_119 (c2670_wire_304, c2670_wire_488_3);
nor_n #(2, 0, 0) NOR_15 (c2670_wire_665, {c2670_wire_666, c2670_wire_302_4});
or_n #(2, 0, 0) OR_95 (c2670_wire_667, {c2670_wire_665, c2670_wire_565});
and_n #(2, 0, 0) AND_240 (c2670_wire_668, {c2670_wire_488_4, c2670_wire_664_1});
or_n #(2, 0, 0) OR_96 (c2670_wire_666, {c2670_wire_668, c2670_wire_305});
notg #(0, 0) NOT_120 (c2670_wire_306, c2670_wire_488_5);
and_n #(2, 0, 0) AND_241 (c2670_wire_669, {c2670_wire_670_0, c2670_wire_488_6});
or_n #(2, 0, 0) OR_97 (c2670_wire_573, {c2670_wire_669, c2670_wire_330});
notg #(0, 0) NOT_121 (c2670_wire_331, c2670_wire_488_7);
nor_n #(2, 0, 0) NOR_16 (c2670_wire_671, {c2670_wire_672, c2670_wire_329_6});
or_n #(2, 0, 0) OR_98 (c2670_wire_673, {c2670_wire_671, c2670_wire_572});
and_n #(2, 0, 0) AND_242 (c2670_wire_674, {c2670_wire_670_1, c2670_wire_488_8});
or_n #(2, 0, 0) OR_99 (c2670_wire_672, {c2670_wire_674, c2670_wire_332});
notg #(0, 0) NOT_122 (c2670_wire_333, c2670_wire_488_9);
and_n #(2, 0, 0) AND_243 (c2670_wire_675, {c2670_wire_676_0, c2670_wire_488_10});
or_n #(2, 0, 0) OR_100 (c2670_wire_600, {c2670_wire_675, c2670_wire_189});
notg #(0, 0) NOT_123 (c2670_wire_190, c2670_wire_488_11);
nor_n #(2, 0, 0) NOR_17 (c2670_wire_677, {c2670_wire_678, c2670_wire_574_4});
or_n #(2, 0, 0) OR_101 (c2670_wire_679, {c2670_wire_677, c2670_wire_599});
and_n #(2, 0, 0) AND_244 (c2670_wire_680, {c2670_wire_676_1, c2670_wire_488_12});
or_n #(2, 0, 0) OR_102 (c2670_wire_678, {c2670_wire_680, c2670_wire_191});
notg #(0, 0) NOT_124 (c2670_wire_192, c2670_wire_488_13);
and_n #(4, 0, 0) AND_245 (c2670_wire_681, {c2670_wire_661, c2670_wire_656, c2670_wire_651, c2670_wire_682});
and_n #(2, 0, 0) AND_246 (c2670_wire_683, {c2670_wire_646, c2670_wire_642});
and_n #(2, 0, 0) AND_247 (c2670_wire_684, {c2670_wire_639, c2670_wire_685});
bufg #(0, 0) BUF_67 (c2670_wire_513, G17_net_0);
and_n #(2, 0, 0) AND_248 (c2670_wire_686, {c2670_wire_679, c2670_wire_673});
and_n #(2, 0, 0) AND_249 (c2670_wire_687, {c2670_wire_667, c2670_wire_688});
and_n #(2, 0, 0) AND_250 (c2670_wire_689, {c2670_wire_276_0, c2670_wire_690});
xor_n #(2, 0, 0) XOR_13 (c2670_wire_690, {c2670_wire_624_0, c2670_wire_626_0});
xor_n #(2, 0, 0) XOR_14 (c2670_wire_691, {c2670_wire_624_1, c2670_wire_626_1});
and_n #(2, 0, 0) AND_251 (c2670_wire_692, {c2670_wire_634_0, c2670_wire_693_0});
and_n #(2, 0, 0) AND_252 (c2670_wire_694, {c2670_wire_634_1, c2670_wire_693_1});
and_n #(2, 0, 0) AND_253 (c2670_wire_682, {c2670_wire_683, c2670_wire_684});
nor_n #(2, 0, 0) NOR_18 (c2670_wire_695, {c2670_wire_110_1, c2670_wire_489_3});
or_n #(2, 0, 0) OR_103 (c2670_wire_696, {c2670_wire_482, c2670_wire_697});
nor_n #(2, 0, 0) NOR_19 (c2670_wire_697, {c2670_wire_371_3, c2670_wire_36_2});
and_n #(3, 0, 0) AND_254 (c2670_wire_698, {c2670_wire_492, c2670_wire_699, c2670_wire_696});
nor_n #(2, 0, 0) NOR_20 (c2670_wire_700, {c2670_wire_489_4, c2670_wire_523_1});
or_n #(2, 0, 0) OR_104 (c2670_wire_494, {c2670_wire_700, c2670_wire_522});
nor_n #(2, 0, 0) NOR_21 (c2670_wire_701, {c2670_wire_371_4, c2670_wire_481_1});
or_n #(2, 0, 0) OR_105 (c2670_wire_495, {c2670_wire_701, c2670_wire_480});
or_n #(2, 0, 0) OR_106 (c2670_wire_699, {c2670_wire_695, c2670_wire_524});
or_n #(2, 0, 0) OR_107 (c2670_wire_685, {c2670_wire_493, c2670_wire_698});
and_n #(2, 0, 0) AND_255 (c2670_wire_702, {c2670_wire_703, c2670_wire_704});
and_n #(2, 0, 0) AND_256 (c2670_wire_703, {c2670_wire_686, c2670_wire_687});
nor_n #(2, 0, 0) NOR_22 (c2670_wire_705, {c2670_wire_347_5, c2670_wire_183_3});
or_n #(2, 0, 0) OR_108 (c2670_wire_706, {c2670_wire_215, c2670_wire_707});
nor_n #(2, 0, 0) NOR_23 (c2670_wire_707, {c2670_wire_209_6, c2670_wire_216_5});
notg #(0, 0) NOT_125 (c2670_wire_708, c2670_wire_488_14);
and_n #(3, 0, 0) AND_257 (c2670_wire_709, {c2670_wire_708, c2670_wire_710, c2670_wire_706});
nor_n #(2, 0, 0) NOR_24 (c2670_wire_711, {c2670_wire_216_6, c2670_wire_602_1});
or_n #(2, 0, 0) OR_109 (c2670_wire_712, {c2670_wire_711, c2670_wire_601});
nor_n #(2, 0, 0) NOR_25 (c2670_wire_713, {c2670_wire_347_6, c2670_wire_577_1});
or_n #(2, 0, 0) OR_110 (c2670_wire_714, {c2670_wire_713, c2670_wire_576});
or_n #(2, 0, 0) OR_111 (c2670_wire_710, {c2670_wire_705, c2670_wire_346});
and_n #(3, 0, 0) AND_258 (c2670_wire_715, {c2670_wire_712, c2670_wire_714, c2670_wire_488_15});
or_n #(2, 0, 0) OR_112 (c2670_wire_688, {c2670_wire_715, c2670_wire_709});
or_n #(2, 0, 0) OR_113 (c2670_wire_716, {c2670_wire_7, c2670_wire_717});
notg #(0, 0) NOT_126 (c2670_wire_718, c2670_wire_716_0);
and_n #(2, 0, 0) AND_259 (c2670_wire_719, {c2670_wire_716_1, c2670_wire_720});
and_n #(2, 0, 0) AND_260 (c2670_wire_721, {c2670_wire_716_2, c2670_wire_722});
nor_n #(2, 0, 0) NOR_26 (c2670_wire_717, {c2670_wire_8_3, c2670_wire_5_7});
bufg #(0, 0) BUF_68 (c2670_wire_518, G18_net_0);
notg #(0, 0) NOT_127 (c2670_wire_723, c2670_wire_386_0);
notg #(0, 0) NOT_128 (c2670_wire_724, c2670_wire_386_1);
or_n #(2, 0, 0) OR_114 (c2670_wire_400, {c2670_wire_618, c2670_wire_725});
or_n #(2, 0, 0) OR_115 (c2670_wire_726, {c2670_wire_620, c2670_wire_727});
or_n #(2, 0, 0) OR_116 (c2670_wire_387, {c2670_wire_399, c2670_wire_728});
nor_n #(2, 0, 0) NOR_27 (c2670_wire_728, {c2670_wire_726, c2670_wire_396_1});
nor_n #(2, 0, 0) NOR_28 (c2670_wire_725, {c2670_wire_585_2, c2670_wire_619_2});
nor_n #(2, 0, 0) NOR_29 (c2670_wire_727, {c2670_wire_585_3, c2670_wire_619_3});
or_n #(2, 0, 0) OR_117 (c2670_wire_405, {c2670_wire_409, c2670_wire_729});
nor_n #(2, 0, 0) NOR_30 (c2670_wire_729, {c2670_wire_406_2, c2670_wire_410_2});
or_n #(2, 0, 0) OR_118 (c2670_wire_730, {c2670_wire_411, c2670_wire_731});
or_n #(2, 0, 0) OR_119 (c2670_wire_732, {c2670_wire_404, c2670_wire_733});
nor_n #(2, 0, 0) NOR_31 (c2670_wire_733, {c2670_wire_730, c2670_wire_401_1});
nor_n #(2, 0, 0) NOR_32 (c2670_wire_731, {c2670_wire_406_3, c2670_wire_410_3});
and_n #(2, 0, 0) AND_261 (c2670_wire_704, {c2670_wire_681, c2670_wire_734});
or_n #(2, 0, 0) OR_120 (c2670_wire_735, {c2670_wire_486, c2670_wire_736});
and_n #(2, 0, 0) AND_262 (c2670_wire_734, {c2670_wire_735, c2670_wire_737});
or_n #(2, 0, 0) OR_121 (c2670_wire_737, {c2670_wire_476, c2670_wire_738});
nor_n #(2, 0, 0) NOR_33 (c2670_wire_736, {c2670_wire_484_1, c2670_wire_284_3});
nor_n #(2, 0, 0) NOR_34 (c2670_wire_738, {c2670_wire_473_1, c2670_wire_477_4});
or_n #(2, 0, 0) OR_122 (c2670_wire_606, {c2670_wire_609, c2670_wire_739});
nor_n #(2, 0, 0) NOR_35 (c2670_wire_739, {c2670_wire_607_3, c2670_wire_610_2});
or_n #(2, 0, 0) OR_123 (c2670_wire_740, {c2670_wire_611, c2670_wire_741});
or_n #(2, 0, 0) OR_124 (c2670_wire_742, {c2670_wire_605, c2670_wire_743});
nor_n #(2, 0, 0) NOR_36 (c2670_wire_743, {c2670_wire_740, c2670_wire_255_2});
nor_n #(2, 0, 0) NOR_37 (c2670_wire_741, {c2670_wire_607_4, c2670_wire_610_3});
notg #(0, 0) NOT_129 (c2670_wire_744, c2670_wire_745);
and_n #(2, 0, 0) AND_263 (c2670_wire_745, {c2670_wire_702, c2670_wire_746});
nor_n #(2, 0, 0) NOR_38 (c2670_wire_747, {c2670_wire_234_5, c2670_wire_604_1});
or_n #(2, 0, 0) OR_125 (c2670_wire_748, {c2670_wire_747, c2670_wire_603});
nor_n #(2, 0, 0) NOR_39 (c2670_wire_749, {c2670_wire_211_4, c2670_wire_234_6});
or_n #(2, 0, 0) OR_126 (c2670_wire_257, {c2670_wire_749, c2670_wire_233});
and_n #(2, 0, 0) AND_264 (c2670_wire_750, {c2670_wire_748, c2670_wire_751});
or_n #(2, 0, 0) OR_127 (c2670_wire_752, {c2670_wire_750, c2670_wire_256});
and_n #(2, 0, 0) AND_265 (c2670_wire_746, {c2670_wire_752, c2670_wire_753});
and_n #(2, 0, 0) AND_266 (c2670_wire_751, {c2670_wire_754, c2670_wire_488_16});
notg #(0, 0) NOT_130 (c2670_wire_258, c2670_wire_488_17);
bufg #(0, 0) BUF_69 (c2670_wire_487, G19_net_0);
and_n #(2, 0, 0) AND_267 (c2670_wire_755, {c2670_wire_756, c2670_wire_757_0});
xor_n #(2, 0, 0) XOR_15 (c2670_wire_758, {c2670_wire_755_0, c2670_wire_759_0});
notg #(0, 0) NOT_131 (c2670_wire_760, c2670_wire_755_1);
notg #(0, 0) NOT_132 (c2670_wire_761, c2670_wire_755_2);
notg #(0, 0) NOT_133 (c2670_wire_756, c2670_wire_110_2);
and_n #(2, 0, 0) AND_268 (c2670_wire_762, {c2670_wire_763, c2670_wire_757_1});
xor_n #(2, 0, 0) XOR_16 (c2670_wire_764, {c2670_wire_762_0, c2670_wire_765_0});
notg #(0, 0) NOT_134 (c2670_wire_766, c2670_wire_762_1);
notg #(0, 0) NOT_135 (c2670_wire_767, c2670_wire_762_2);
notg #(0, 0) NOT_136 (c2670_wire_763, c2670_wire_126_2);
and_n #(2, 0, 0) AND_269 (c2670_wire_768, {c2670_wire_34_0, c2670_wire_612});
xor_n #(2, 0, 0) XOR_17 (c2670_wire_722, {c2670_wire_34_1, c2670_wire_769_0});
xor_n #(2, 0, 0) XOR_18 (c2670_wire_770, {c2670_wire_34_2, c2670_wire_769_1});
xor_n #(2, 0, 0) XOR_19 (c2670_wire_769, {c2670_wire_91_3, c2670_wire_110_3});
or_n #(2, 0, 0) OR_128 (c2670_wire_771, {c2670_wire_772, c2670_wire_773});
and_n #(2, 0, 0) AND_270 (c2670_wire_774, {c2670_wire_771_0, c2670_wire_775});
and_n #(2, 0, 0) AND_271 (c2670_wire_772, {c2670_wire_157_1, c2670_wire_173_3});
nor_n #(2, 0, 0) NOR_40 (c2670_wire_773, {c2670_wire_157_2, c2670_wire_173_4});
and_n #(2, 0, 0) AND_272 (c2670_wire_776, {c2670_wire_11, c2670_wire_40});
and_n #(2, 0, 0) AND_273 (c2670_wire_777, {c2670_wire_12, c2670_wire_39});
or_n #(2, 0, 0) OR_129 (c2670_wire_452, {c2670_wire_777, c2670_wire_776});
bufg #(0, 0) BUF_70 (c2670_wire_440, G2_net_0);
bufg #(0, 0) BUF_71 (c2670_wire_670, G20_net_0);
nor_n #(2, 0, 0) NOR_41 (c2670_wire_778, {c2670_wire_276_1, c2670_wire_691});
or_n #(2, 0, 0) OR_130 (c2670_wire_693, {c2670_wire_689, c2670_wire_778});
bufg #(0, 0) BUF_72 (c2670_wire_676, G21_net_0);
or_n #(2, 0, 0) OR_131 (c2670_wire_779, {c2670_wire_528, c2670_wire_780});
and_n #(2, 0, 0) AND_274 (c2670_wire_781, {c2670_wire_779_0, c2670_wire_782_0});
or_n #(2, 0, 0) OR_132 (c2670_wire_783, {c2670_wire_779_1, c2670_wire_782_1});
and_n #(2, 0, 0) AND_275 (c2670_wire_784, {c2670_wire_779_2, c2670_wire_782_2});
or_n #(2, 0, 0) OR_133 (c2670_wire_785, {c2670_wire_779_3, c2670_wire_782_3});
nor_n #(2, 0, 0) NOR_42 (c2670_wire_780, {c2670_wire_466_3, c2670_wire_526_16});
and_n #(2, 0, 0) AND_276 (c2670_wire_786, {c2670_wire_787_0, c2670_wire_36_3});
or_n #(2, 0, 0) OR_134 (c2670_wire_787, {c2670_wire_530, c2670_wire_788});
and_n #(2, 0, 0) AND_277 (c2670_wire_789, {c2670_wire_787_1, c2670_wire_36_4});
and_n #(2, 0, 0) AND_278 (c2670_wire_790, {c2670_wire_787_2, c2670_wire_36_5});
nor_n #(2, 0, 0) NOR_43 (c2670_wire_788, {c2670_wire_371_5, c2670_wire_526_17});
and_n #(2, 0, 0) AND_279 (c2670_wire_791, {c2670_wire_792_0, c2670_wire_91_4});
or_n #(2, 0, 0) OR_135 (c2670_wire_792, {c2670_wire_532, c2670_wire_793});
and_n #(2, 0, 0) AND_280 (c2670_wire_794, {c2670_wire_792_1, c2670_wire_91_5});
and_n #(2, 0, 0) AND_281 (c2670_wire_795, {c2670_wire_792_2, c2670_wire_91_6});
nor_n #(2, 0, 0) NOR_44 (c2670_wire_793, {c2670_wire_483_3, c2670_wire_526_18});
bufg #(0, 0) BUF_73 (c2670_wire_754, G22_net_0);
and_n #(2, 0, 0) AND_282 (c2670_wire_796, {c2670_wire_718, c2670_wire_797});
or_n #(2, 0, 0) OR_136 (c2670_wire_798, {c2670_wire_796_0, c2670_wire_719_0});
notg #(0, 0) NOT_137 (c2670_wire_799, c2670_wire_796_1);
and_n #(3, 0, 0) AND_283 (c2670_wire_800, {c2670_wire_432, c2670_wire_42, c2670_wire_36_6});
nor_n #(2, 0, 0) NOR_45 (c2670_wire_801, {c2670_wire_459_2, c2670_wire_34_3});
or_n #(2, 0, 0) OR_137 (c2670_wire_797, {c2670_wire_800, c2670_wire_801});
notg #(0, 0) NOT_138 (c2670_wire_802, c2670_wire_719_1);
nor_n #(3, 0, 0) NOR_46 (c2670_wire_803, {c2670_wire_13_5, c2670_wire_35_10, c2670_wire_36_7});
or_n #(2, 0, 0) OR_138 (c2670_wire_720, {c2670_wire_768, c2670_wire_803});
and_n #(2, 0, 0) AND_284 (c2670_wire_804, {c2670_wire_805_0, c2670_wire_806_0});
notg #(0, 0) NOT_139 (c2670_wire_807, c2670_wire_805_1);
and_n #(3, 0, 0) AND_285 (c2670_wire_808, {c2670_wire_805_2, c2670_wire_802, c2670_wire_799});
or_n #(2, 0, 0) OR_139 (c2670_wire_805, {c2670_wire_774, c2670_wire_809});
and_n #(2, 0, 0) AND_286 (c2670_wire_810, {c2670_wire_126_3, c2670_wire_147_2});
or_n #(2, 0, 0) OR_140 (c2670_wire_775, {c2670_wire_810, c2670_wire_811});
or_n #(2, 0, 0) OR_141 (c2670_wire_812, {c2670_wire_813, c2670_wire_814});
nor_n #(2, 0, 0) NOR_47 (c2670_wire_809, {c2670_wire_812, c2670_wire_771_1});
nor_n #(2, 0, 0) NOR_48 (c2670_wire_811, {c2670_wire_126_4, c2670_wire_147_3});
and_n #(2, 0, 0) AND_287 (c2670_wire_813, {c2670_wire_126_5, c2670_wire_147_4});
nor_n #(2, 0, 0) NOR_49 (c2670_wire_814, {c2670_wire_126_6, c2670_wire_147_5});
and_n #(2, 0, 0) AND_288 (c2670_wire_782, {c2670_wire_14, c2670_wire_815});
nor_n #(2, 0, 0) NOR_50 (c2670_wire_816, {c2670_wire_465_3, c2670_wire_526_19});
or_n #(2, 0, 0) OR_142 (c2670_wire_815, {c2670_wire_536, c2670_wire_816});
and_n #(2, 0, 0) AND_289 (c2670_wire_759, {c2670_wire_817, c2670_wire_757_2});
and_n #(2, 0, 0) AND_290 (c2670_wire_818, {c2670_wire_759_1, c2670_wire_760});
and_n #(2, 0, 0) AND_291 (c2670_wire_819, {c2670_wire_759_2, c2670_wire_761});
nor_n #(2, 0, 0) NOR_51 (c2670_wire_820, {c2670_wire_489_5, c2670_wire_526_20});
or_n #(2, 0, 0) OR_143 (c2670_wire_817, {c2670_wire_538, c2670_wire_820});
and_n #(2, 0, 0) AND_292 (c2670_wire_765, {c2670_wire_821, c2670_wire_757_3});
and_n #(2, 0, 0) AND_293 (c2670_wire_822, {c2670_wire_765_1, c2670_wire_766});
and_n #(2, 0, 0) AND_294 (c2670_wire_823, {c2670_wire_765_2, c2670_wire_767});
nor_n #(2, 0, 0) NOR_52 (c2670_wire_824, {c2670_wire_525_3, c2670_wire_526_21});
or_n #(2, 0, 0) OR_144 (c2670_wire_821, {c2670_wire_534, c2670_wire_824});
nor_n #(2, 0, 0) NOR_53 (c2670_wire_825, {c2670_wire_716_3, c2670_wire_770});
or_n #(2, 0, 0) OR_145 (c2670_wire_806, {c2670_wire_721, c2670_wire_825});
bufg #(0, 0) BUF_74 (c2670_wire_488, G23_net_0);
notg #(0, 0) NOT_140 (c2670_wire_826, c2670_wire_827_0);
notg #(0, 0) NOT_141 (c2670_wire_828, c2670_wire_827_1);
and_n #(2, 0, 0) AND_295 (c2670_wire_827, {c2670_wire_829, c2670_wire_830});
or_n #(2, 0, 0) OR_146 (c2670_wire_260, {c2670_wire_692, c2670_wire_831});
nor_n #(2, 0, 0) NOR_54 (c2670_wire_832, {c2670_wire_634_2, c2670_wire_693_2});
or_n #(2, 0, 0) OR_147 (c2670_wire_833, {c2670_wire_832, c2670_wire_694});
or_n #(2, 0, 0) OR_148 (c2670_wire_829, {c2670_wire_259, c2670_wire_834});
nor_n #(2, 0, 0) NOR_55 (c2670_wire_834, {c2670_wire_833, c2670_wire_251_3});
nor_n #(2, 0, 0) NOR_56 (c2670_wire_831, {c2670_wire_634_3, c2670_wire_693_3});
notg #(0, 0) NOT_142 (c2670_wire_830, c2670_wire_835_0);
notg #(0, 0) NOT_143 (c2670_wire_836, c2670_wire_596_0);
notg #(0, 0) NOT_144 (c2670_wire_837, c2670_wire_596_1);
notg #(0, 0) NOT_145 (c2670_wire_838, c2670_wire_594_0);
notg #(0, 0) NOT_146 (c2670_wire_839, c2670_wire_594_1);
or_n #(2, 0, 0) OR_149 (c2670_wire_595, {c2670_wire_301, c2670_wire_840});
nor_n #(2, 0, 0) NOR_57 (c2670_wire_840, {c2670_wire_297_5, c2670_wire_302_5});
notg #(0, 0) NOT_147 (c2670_wire_841, c2670_wire_597_0);
notg #(0, 0) NOT_148 (c2670_wire_842, c2670_wire_597_1);
or_n #(2, 0, 0) OR_150 (c2670_wire_598, {c2670_wire_283, c2670_wire_843});
nor_n #(2, 0, 0) NOR_58 (c2670_wire_843, {c2670_wire_277_3, c2670_wire_284_4});
notg #(0, 0) NOT_149 (c2670_wire_844, c2670_wire_593_0);
notg #(0, 0) NOT_150 (c2670_wire_845, c2670_wire_846_0);
and_n #(2, 0, 0) AND_296 (c2670_wire_846, {c2670_wire_847, c2670_wire_757_4});
notg #(0, 0) NOT_151 (c2670_wire_547, c2670_wire_157_3);
nor_n #(2, 0, 0) NOR_59 (c2670_wire_848, {c2670_wire_526_22, c2670_wire_477_5});
or_n #(2, 0, 0) OR_151 (c2670_wire_847, {c2670_wire_546, c2670_wire_848});
notg #(0, 0) NOT_152 (c2670_wire_849, c2670_wire_850_0);
notg #(0, 0) NOT_153 (c2670_wire_851, c2670_wire_850_1);
and_n #(2, 0, 0) AND_297 (c2670_wire_850, {c2670_wire_852, c2670_wire_757_5});
notg #(0, 0) NOT_154 (c2670_wire_545, c2670_wire_147_6);
nor_n #(2, 0, 0) NOR_60 (c2670_wire_853, {c2670_wire_526_23, c2670_wire_552_3});
or_n #(2, 0, 0) OR_152 (c2670_wire_852, {c2670_wire_544, c2670_wire_853});
bufg #(0, 0) BUF_75 (c2670_wire_664, G24_net_0);
or_n #(2, 0, 0) OR_153 (c2670_wire_854, {c2670_wire_786, c2670_wire_855});
notg #(0, 0) NOT_155 (c2670_wire_856, c2670_wire_854_0);
notg #(0, 0) NOT_156 (c2670_wire_857, c2670_wire_854_1);
nor_n #(2, 0, 0) NOR_61 (c2670_wire_855, {c2670_wire_36_8, c2670_wire_787_3});
or_n #(2, 0, 0) OR_154 (c2670_wire_858, {c2670_wire_791, c2670_wire_859});
notg #(0, 0) NOT_157 (c2670_wire_860, c2670_wire_858_0);
notg #(0, 0) NOT_158 (c2670_wire_861, c2670_wire_858_1);
nor_n #(2, 0, 0) NOR_62 (c2670_wire_859, {c2670_wire_91_7, c2670_wire_792_3});
nor_n #(4, 0, 0) NOR_63 (c2670_wire_862, {c2670_wire_594_2, c2670_wire_593_1, c2670_wire_597_2, c2670_wire_596_2});
and_n #(2, 0, 0) AND_298 (c2670_wire_863, {c2670_wire_862_0, c2670_wire_864_0});
notg #(0, 0) NOT_159 (c2670_wire_865, c2670_wire_764_0);
notg #(0, 0) NOT_160 (c2670_wire_866, c2670_wire_764_1);
notg #(0, 0) NOT_161 (c2670_wire_867, c2670_wire_758_0);
notg #(0, 0) NOT_162 (c2670_wire_868, c2670_wire_758_1);
notg #(0, 0) NOT_163 (c2670_wire_869, c2670_wire_587_0);
or_n #(2, 0, 0) OR_155 (c2670_wire_870, {c2670_wire_587_1, c2670_wire_863});
or_n #(2, 0, 0) OR_156 (c2670_wire_588, {c2670_wire_324, c2670_wire_871});
and_n #(3, 0, 0) AND_299 (c2670_wire_872, {c2670_wire_841, c2670_wire_560, c2670_wire_173_5});
or_n #(2, 0, 0) OR_157 (c2670_wire_873, {c2670_wire_872, c2670_wire_874});
nor_n #(2, 0, 0) NOR_64 (c2670_wire_874, {c2670_wire_277_4, c2670_wire_284_5});
nor_n #(2, 0, 0) NOR_65 (c2670_wire_875, {c2670_wire_297_6, c2670_wire_302_6});
or_n #(2, 0, 0) OR_158 (c2670_wire_876, {c2670_wire_875, c2670_wire_877});
and_n #(2, 0, 0) AND_300 (c2670_wire_877, {c2670_wire_873, c2670_wire_838});
and_n #(2, 0, 0) AND_301 (c2670_wire_871, {c2670_wire_876, c2670_wire_836});
notg #(0, 0) NOT_164 (c2670_wire_878, c2670_wire_879_0);
and_n #(2, 0, 0) AND_302 (c2670_wire_879, {c2670_wire_880, c2670_wire_881});
notg #(0, 0) NOT_165 (c2670_wire_882, c2670_wire_879_1);
or_n #(2, 0, 0) OR_159 (c2670_wire_881, {c2670_wire_804, c2670_wire_883});
nor_n #(2, 0, 0) NOR_66 (c2670_wire_883, {c2670_wire_805_3, c2670_wire_806_1});
notg #(0, 0) NOT_166 (c2670_wire_880, c2670_wire_835_1);
or_n #(2, 0, 0) OR_160 (c2670_wire_864, {c2670_wire_884, c2670_wire_885});
nor_n #(2, 0, 0) NOR_67 (c2670_wire_886, {c2670_wire_552_4, c2670_wire_846_1});
and_n #(2, 0, 0) AND_303 (c2670_wire_887, {c2670_wire_783, c2670_wire_43});
and_n #(2, 0, 0) AND_304 (c2670_wire_888, {c2670_wire_856, c2670_wire_889});
and_n #(2, 0, 0) AND_305 (c2670_wire_890, {c2670_wire_860, c2670_wire_891});
and_n #(2, 0, 0) AND_306 (c2670_wire_892, {c2670_wire_867, c2670_wire_893});
and_n #(2, 0, 0) AND_307 (c2670_wire_894, {c2670_wire_865, c2670_wire_895});
and_n #(3, 0, 0) AND_308 (c2670_wire_885, {c2670_wire_849, c2670_wire_845, c2670_wire_896});
or_n #(2, 0, 0) OR_161 (c2670_wire_897, {c2670_wire_886, c2670_wire_558});
or_n #(2, 0, 0) OR_162 (c2670_wire_896, {c2670_wire_822, c2670_wire_894});
or_n #(2, 0, 0) OR_163 (c2670_wire_895, {c2670_wire_818, c2670_wire_892});
or_n #(2, 0, 0) OR_164 (c2670_wire_889, {c2670_wire_887, c2670_wire_781});
and_n #(3, 0, 0) AND_309 (c2670_wire_884, {c2670_wire_897, c2670_wire_541, c2670_wire_757_6});
or_n #(2, 0, 0) OR_165 (c2670_wire_891, {c2670_wire_888, c2670_wire_789});
or_n #(2, 0, 0) OR_166 (c2670_wire_893, {c2670_wire_890, c2670_wire_794});
bufg #(0, 0) BUF_76 (c2670_wire_577, G25_net_0);
notg #(0, 0) NOT_167 (c2670_wire_898, c2670_wire_899_0);
notg #(0, 0) NOT_168 (c2670_wire_900, c2670_wire_899_1);
and_n #(3, 0, 0) AND_310 (c2670_wire_901, {c2670_wire_899_2, c2670_wire_869, c2670_wire_902});
or_n #(2, 0, 0) OR_167 (c2670_wire_899, {c2670_wire_589, c2670_wire_903});
nor_n #(2, 0, 0) NOR_68 (c2670_wire_904, {c2670_wire_552_5, c2670_wire_846_2});
or_n #(2, 0, 0) OR_168 (c2670_wire_905, {c2670_wire_559, c2670_wire_904});
nor_n #(2, 0, 0) NOR_69 (c2670_wire_906, {c2670_wire_597_3, c2670_wire_593_2});
and_n #(2, 0, 0) AND_311 (c2670_wire_907, {c2670_wire_543, c2670_wire_908});
or_n #(2, 0, 0) OR_169 (c2670_wire_909, {c2670_wire_795, c2670_wire_910});
or_n #(2, 0, 0) OR_170 (c2670_wire_911, {c2670_wire_790, c2670_wire_912});
nor_n #(3, 0, 0) NOR_70 (c2670_wire_913, {c2670_wire_302_7, c2670_wire_297_7, c2670_wire_596_3});
or_n #(2, 0, 0) OR_171 (c2670_wire_914, {c2670_wire_784, c2670_wire_915});
and_n #(2, 0, 0) AND_312 (c2670_wire_915, {c2670_wire_785, c2670_wire_44});
and_n #(2, 0, 0) AND_313 (c2670_wire_912, {c2670_wire_857, c2670_wire_914});
and_n #(2, 0, 0) AND_314 (c2670_wire_910, {c2670_wire_861, c2670_wire_911});
and_n #(2, 0, 0) AND_315 (c2670_wire_916, {c2670_wire_868, c2670_wire_909});
and_n #(2, 0, 0) AND_316 (c2670_wire_917, {c2670_wire_866, c2670_wire_918});
and_n #(3, 0, 0) AND_317 (c2670_wire_919, {c2670_wire_844, c2670_wire_920, c2670_wire_921});
nor_n #(2, 0, 0) NOR_71 (c2670_wire_920, {c2670_wire_597_4, c2670_wire_846_3});
and_n #(2, 0, 0) AND_318 (c2670_wire_922, {c2670_wire_851, c2670_wire_919});
and_n #(3, 0, 0) AND_319 (c2670_wire_903, {c2670_wire_839, c2670_wire_837, c2670_wire_923});
or_n #(2, 0, 0) OR_172 (c2670_wire_590, {c2670_wire_326, c2670_wire_913});
and_n #(3, 0, 0) AND_320 (c2670_wire_924, {c2670_wire_842, c2670_wire_561, c2670_wire_173_6});
or_n #(2, 0, 0) OR_173 (c2670_wire_592, {c2670_wire_924, c2670_wire_925});
nor_n #(2, 0, 0) NOR_72 (c2670_wire_925, {c2670_wire_277_5, c2670_wire_284_6});
and_n #(3, 0, 0) AND_321 (c2670_wire_926, {c2670_wire_906, c2670_wire_905, c2670_wire_757_7});
or_n #(2, 0, 0) OR_174 (c2670_wire_921, {c2670_wire_823, c2670_wire_917});
or_n #(2, 0, 0) OR_175 (c2670_wire_918, {c2670_wire_819, c2670_wire_916});
or_n #(2, 0, 0) OR_176 (c2670_wire_908, {c2670_wire_591, c2670_wire_926});
or_n #(2, 0, 0) OR_177 (c2670_wire_923, {c2670_wire_907, c2670_wire_922});
and_n #(2, 0, 0) AND_322 (c2670_wire_927, {c2670_wire_900, c2670_wire_870});
nand_n #(2, 0, 0) NAND_2 (c2670_wire_902, {c2670_wire_862_1, c2670_wire_864_1});
or_n #(2, 0, 0) OR_178 (c2670_wire_928, {c2670_wire_927, c2670_wire_901});
notg #(0, 0) NOT_169 (c2670_wire_929, c2670_wire_930);
and_n #(7, 0, 0) AND_323 (c2670_wire_930, {c2670_wire_828, c2670_wire_882, c2670_wire_931, c2670_wire_724, c2670_wire_932, c2670_wire_933, c2670_wire_420_2});
notg #(0, 0) NOT_170 (c2670_wire_931, c2670_wire_742_0);
notg #(0, 0) NOT_171 (c2670_wire_932, c2670_wire_732_0);
notg #(0, 0) NOT_172 (c2670_wire_933, c2670_wire_928_0);
bufg #(0, 0) BUF_77 (G2531_net_0, c2670_wire_934_0);
bufg #(0, 0) BUF_78 (G2532_net_0, c2670_wire_934_1);
notg #(0, 0) NOT_173 (c2670_wire_934, c2670_wire_428_0);
bufg #(0, 0) BUF_79 (G2533_net_0, c2670_wire_934_2);
bufg #(0, 0) BUF_80 (G2534_net_0, c2670_wire_464_0);
bufg #(0, 0) BUF_81 (G2535_net_0, c2670_wire_464_1);
bufg #(0, 0) BUF_82 (G2536_net_0, c2670_wire_571_0);
bufg #(0, 0) BUF_83 (G2537_net_0, c2670_wire_571_1);
bufg #(0, 0) BUF_84 (G2538_net_0, c2670_wire_571_2);
bufg #(0, 0) BUF_85 (G2539_net_0, c2670_wire_935);
notg #(0, 0) NOT_174 (c2670_wire_935, c2670_wire_319_1);
bufg #(0, 0) BUF_86 (G2540_net_0, c2670_wire_317);
bufg #(0, 0) BUF_87 (G2541_net_0, c2670_wire_936);
notg #(0, 0) NOT_175 (c2670_wire_936, c2670_wire_320_1);
bufg #(0, 0) BUF_88 (G2542_net_0, c2670_wire_937);
notg #(0, 0) NOT_176 (c2670_wire_937, c2670_wire_321_1);
bufg #(0, 0) BUF_89 (G2543_net_0, c2670_wire_938);
notg #(0, 0) NOT_177 (c2670_wire_938, c2670_wire_939_0);
bufg #(0, 0) BUF_90 (G2544_net_0, c2670_wire_940);
notg #(0, 0) NOT_178 (c2670_wire_940, c2670_wire_941_0);
bufg #(0, 0) BUF_91 (G2545_net_0, c2670_wire_942);
notg #(0, 0) NOT_179 (c2670_wire_942, c2670_wire_943_0);
bufg #(0, 0) BUF_92 (G2546_net_0, c2670_wire_944);
notg #(0, 0) NOT_180 (c2670_wire_944, c2670_wire_945_0);
bufg #(0, 0) BUF_93 (G2547_net_0, c2670_wire_946);
notg #(0, 0) NOT_181 (c2670_wire_946, c2670_wire_575);
bufg #(0, 0) BUF_94 (G2548_net_0, c2670_wire_947);
notg #(0, 0) NOT_182 (c2670_wire_947, c2670_wire_439);
bufg #(0, 0) BUF_95 (G2549_net_0, c2670_wire_428_1);
notg #(0, 0) NOT_183 (c2670_wire_948, c2670_wire_428_2);
bufg #(0, 0) BUF_96 (G2550_net_0, c2670_wire_949);
and_n #(2, 0, 0) AND_324 (c2670_wire_949, {c2670_wire_948, c2670_wire_950});
bufg #(0, 0) BUF_97 (G2551_net_0, c2670_wire_951);
nand_n #(2, 0, 0) NAND_3 (c2670_wire_951, {c2670_wire_419_5, c2670_wire_438_2});
bufg #(0, 0) BUF_98 (G2552_net_0, c2670_wire_952);
notg #(0, 0) NOT_184 (c2670_wire_952, c2670_wire_437);
bufg #(0, 0) BUF_99 (G2553_net_0, c2670_wire_953);
notg #(0, 0) NOT_185 (c2670_wire_953, c2670_wire_448);
bufg #(0, 0) BUF_100 (G2554_net_0, c2670_wire_954_0);
bufg #(0, 0) BUF_101 (G2555_net_0, c2670_wire_954_1);
nand_n #(2, 0, 0) NAND_4 (c2670_wire_954, {c2670_wire_318_0, c2670_wire_955_0});
bufg #(0, 0) BUF_102 (G2556_net_0, c2670_wire_956);
notg #(0, 0) NOT_186 (c2670_wire_956, c2670_wire_420_3);
bufg #(0, 0) BUF_103 (G2557_net_0, c2670_wire_208);
bufg #(0, 0) BUF_104 (G2558_net_0, c2670_wire_230);
bufg #(0, 0) BUF_105 (G2559_net_0, c2670_wire_180);
bufg #(0, 0) BUF_106 (G2560_net_0, c2670_wire_957);
notg #(0, 0) NOT_187 (c2670_wire_957, c2670_wire_126_7);
bufg #(0, 0) BUF_107 (G2561_net_0, c2670_wire_958);
notg #(0, 0) NOT_188 (c2670_wire_958, c2670_wire_110_4);
bufg #(0, 0) BUF_108 (G2562_net_0, c2670_wire_959);
notg #(0, 0) NOT_189 (c2670_wire_959, c2670_wire_91_8);
bufg #(0, 0) BUF_109 (G2563_net_0, c2670_wire_4);
bufg #(0, 0) BUF_110 (G2564_net_0, c2670_wire_412);
bufg #(0, 0) BUF_111 (G2565_net_0, c2670_wire_421);
bufg #(0, 0) BUF_112 (G2566_net_0, c2670_wire_36_9);
and_n #(2, 0, 0) AND_325 (c2670_wire_960, {c2670_wire_36_10, c2670_wire_454});
bufg #(0, 0) BUF_113 (G2567_net_0, c2670_wire_91_9);
bufg #(0, 0) BUF_114 (G2568_net_0, c2670_wire_110_5);
notg #(0, 0) NOT_190 (c2670_wire_456, c2670_wire_110_6);
bufg #(0, 0) BUF_115 (G2569_net_0, c2670_wire_126_8);
bufg #(0, 0) BUF_116 (G2570_net_0, c2670_wire_147_7);
bufg #(0, 0) BUF_117 (G2571_net_0, c2670_wire_157_4);
bufg #(0, 0) BUF_118 (G2572_net_0, c2670_wire_173_7);
bufg #(0, 0) BUF_119 (G2573_net_0, c2670_wire_961_0);
bufg #(0, 0) BUF_120 (G2574_net_0, c2670_wire_961_1);
or_n #(2, 0, 0) OR_179 (c2670_wire_961, {c2670_wire_457, c2670_wire_962});
nor_n #(2, 0, 0) NOR_73 (c2670_wire_962, {c2670_wire_453_6, c2670_wire_35_11});
bufg #(0, 0) BUF_121 (G2575_net_0, c2670_wire_963_0);
bufg #(0, 0) BUF_122 (G2576_net_0, c2670_wire_963_1);
or_n #(2, 0, 0) OR_180 (c2670_wire_963, {c2670_wire_960, c2670_wire_455});
bufg #(0, 0) BUF_123 (G2577_net_0, c2670_wire_49);
bufg #(0, 0) BUF_124 (G2578_net_0, c2670_wire_964_0);
bufg #(0, 0) BUF_125 (G2579_net_0, c2670_wire_964_1);
or_n #(2, 0, 0) OR_181 (c2670_wire_964, {c2670_wire_458, c2670_wire_965});
nor_n #(2, 0, 0) NOR_74 (c2670_wire_965, {c2670_wire_453_7, c2670_wire_5_8});
bufg #(0, 0) BUF_126 (G2580_net_0, c2670_wire_966);
nor_n #(2, 0, 0) NOR_75 (c2670_wire_967, {c2670_wire_255_3, c2670_wire_251_4});
or_n #(2, 0, 0) OR_182 (c2670_wire_966, {c2670_wire_608, c2670_wire_967});
bufg #(0, 0) BUF_127 (G2581_net_0, c2670_wire_723);
bufg #(0, 0) BUF_128 (G2582_net_0, c2670_wire_742_1);
bufg #(0, 0) BUF_129 (G2583_net_0, c2670_wire_732_1);
bufg #(0, 0) BUF_130 (G2584_net_0, c2670_wire_744_0);
bufg #(0, 0) BUF_131 (G2585_net_0, c2670_wire_744_1);
bufg #(0, 0) BUF_132 (G2586_net_0, c2670_wire_968);
nor_n #(3, 0, 0) NOR_76 (c2670_wire_969, {c2670_wire_8_4, c2670_wire_450_3, c2670_wire_452_1});
or_n #(2, 0, 0) OR_183 (c2670_wire_968, {c2670_wire_569, c2670_wire_969});
bufg #(0, 0) BUF_133 (G2587_net_0, c2670_wire_826);
bufg #(0, 0) BUF_134 (G2588_net_0, c2670_wire_970_0);
bufg #(0, 0) BUF_135 (G2589_net_0, c2670_wire_970_1);
and_n #(2, 0, 0) AND_326 (c2670_wire_971, {c2670_wire_798, c2670_wire_807});
or_n #(2, 0, 0) OR_184 (c2670_wire_970, {c2670_wire_461, c2670_wire_570});
or_n #(2, 0, 0) OR_185 (c2670_wire_462, {c2670_wire_971, c2670_wire_808});
bufg #(0, 0) BUF_136 (G2590_net_0, c2670_wire_878);
bufg #(0, 0) BUF_137 (G2591_net_0, c2670_wire_898);
bufg #(0, 0) BUF_138 (G2592_net_0, c2670_wire_928_1);
bufg #(0, 0) BUF_139 (G2593_net_0, c2670_wire_929_0);
bufg #(0, 0) BUF_140 (G2594_net_0, c2670_wire_929_1);
bufg #(0, 0) BUF_141 (c2670_wire_602, G26_net_0);
bufg #(0, 0) BUF_142 (c2670_wire_604, G27_net_0);
bufg #(0, 0) BUF_143 (c2670_wire_417, G28_net_0);
bufg #(0, 0) BUF_144 (c2670_wire_835, G29_net_0);
bufg #(0, 0) BUF_145 (c2670_wire_426, G3_net_0);
bufg #(0, 0) BUF_146 (c2670_wire_187, G30_net_0);
bufg #(0, 0) BUF_147 (c2670_wire_30, G31_net_0);
bufg #(0, 0) BUF_148 (c2670_wire_319, G32_net_0);
bufg #(0, 0) BUF_149 (c2670_wire_176, G33_net_0);
or_n #(2, 0, 0) OR_186 (c2670_wire_972, {c2670_wire_318_1, c2670_wire_613});
notg #(0, 0) NOT_191 (c2670_wire_436, c2670_wire_955_1);
and_n #(4, 0, 0) AND_327 (c2670_wire_955, {c2670_wire_943_1, c2670_wire_939_1, c2670_wire_945_1, c2670_wire_941_1});
bufg #(0, 0) BUF_150 (c2670_wire_160, G34_net_0);
bufg #(0, 0) BUF_151 (c2670_wire_143, G35_net_0);
bufg #(0, 0) BUF_152 (c2670_wire_129, G36_net_0);
bufg #(0, 0) BUF_153 (c2670_wire_113, G37_net_0);
bufg #(0, 0) BUF_154 (c2670_wire_94, G38_net_0);
bufg #(0, 0) BUF_155 (c2670_wire_78, G39_net_0);
bufg #(0, 0) BUF_156 (c2670_wire_510, G4_net_0);
bufg #(0, 0) BUF_157 (c2670_wire_60, G40_net_0);
bufg #(0, 0) BUF_158 (c2670_wire_446, G41_net_0);
bufg #(0, 0) BUF_159 (c2670_wire_28, G42_net_0);
bufg #(0, 0) BUF_160 (c2670_wire_943, G43_net_0);
bufg #(0, 0) BUF_161 (c2670_wire_169, G44_net_0);
bufg #(0, 0) BUF_162 (c2670_wire_153, G45_net_0);
bufg #(0, 0) BUF_163 (c2670_wire_122, G46_net_0);
bufg #(0, 0) BUF_164 (c2670_wire_106, G47_net_0);
bufg #(0, 0) BUF_165 (c2670_wire_87, G48_net_0);
bufg #(0, 0) BUF_166 (c2670_wire_72, G49_net_0);
bufg #(0, 0) BUF_167 (c2670_wire_500, G5_net_0);
bufg #(0, 0) BUF_168 (c2670_wire_58, G50_net_0);
bufg #(0, 0) BUF_169 (c2670_wire_973, G51_net_0);
and_n #(2, 0, 0) AND_328 (c2670_wire_974, {c2670_wire_973, c2670_wire_444});
bufg #(0, 0) BUF_170 (c2670_wire_33, G52_net_0);
bufg #(0, 0) BUF_171 (c2670_wire_939, G53_net_0);
bufg #(0, 0) BUF_172 (c2670_wire_179, G54_net_0);
bufg #(0, 0) BUF_173 (c2670_wire_163, G55_net_0);
bufg #(0, 0) BUF_174 (c2670_wire_141, G56_net_0);
bufg #(0, 0) BUF_175 (c2670_wire_132, G57_net_0);
bufg #(0, 0) BUF_176 (c2670_wire_116, G58_net_0);
bufg #(0, 0) BUF_177 (c2670_wire_97, G59_net_0);
bufg #(0, 0) BUF_178 (c2670_wire_478, G6_net_0);
bufg #(0, 0) BUF_179 (c2670_wire_81, G60_net_0);
bufg #(0, 0) BUF_180 (c2670_wire_63, G61_net_0);
bufg #(0, 0) BUF_181 (c2670_wire_975, G62_net_0);
and_n #(2, 0, 0) AND_329 (c2670_wire_976, {c2670_wire_975, c2670_wire_447});
bufg #(0, 0) BUF_182 (c2670_wire_21, G63_net_0);
bufg #(0, 0) BUF_183 (c2670_wire_320, G64_net_0);
bufg #(0, 0) BUF_184 (c2670_wire_165, G65_net_0);
bufg #(0, 0) BUF_185 (c2670_wire_149, G66_net_0);
bufg #(0, 0) BUF_186 (c2670_wire_138, G67_net_0);
bufg #(0, 0) BUF_187 (c2670_wire_118, G68_net_0);
bufg #(0, 0) BUF_188 (c2670_wire_102, G69_net_0);
or_n #(2, 0, 0) OR_187 (c2670_wire_582, {c2670_wire_615, c2670_wire_977});
nor_n #(2, 0, 0) NOR_77 (c2670_wire_977, {c2670_wire_616_1, c2670_wire_614_1});
or_n #(2, 0, 0) OR_188 (c2670_wire_579, {c2670_wire_621, c2670_wire_978});
nor_n #(2, 0, 0) NOR_78 (c2670_wire_978, {c2670_wire_622_1, c2670_wire_617_1});
or_n #(2, 0, 0) OR_189 (c2670_wire_580, {c2670_wire_628, c2670_wire_979});
nor_n #(2, 0, 0) NOR_79 (c2670_wire_979, {c2670_wire_629_1, c2670_wire_623_1});
bufg #(0, 0) BUF_189 (c2670_wire_438, G7_net_0);
bufg #(0, 0) BUF_190 (c2670_wire_83, G70_net_0);
bufg #(0, 0) BUF_191 (c2670_wire_68, G71_net_0);
bufg #(0, 0) BUF_192 (c2670_wire_52, G72_net_0);
bufg #(0, 0) BUF_193 (c2670_wire_443, G73_net_0);
bufg #(0, 0) BUF_194 (c2670_wire_950, G74_net_0);
bufg #(0, 0) BUF_195 (c2670_wire_292, G75_net_0);
bufg #(0, 0) BUF_196 (c2670_wire_321, G76_net_0);
bufg #(0, 0) BUF_197 (c2670_wire_270, G77_net_0);
or_n #(2, 0, 0) OR_190 (c2670_wire_619, {c2670_wire_631, c2670_wire_980});
nor_n #(2, 0, 0) NOR_80 (c2670_wire_980, {c2670_wire_632_1, c2670_wire_630_1});
bufg #(0, 0) BUF_198 (c2670_wire_244, G78_net_0);
bufg #(0, 0) BUF_199 (c2670_wire_226, G79_net_0);
bufg #(0, 0) BUF_200 (c2670_wire_757, G8_net_0);
bufg #(0, 0) BUF_201 (c2670_wire_201, G80_net_0);
bufg #(0, 0) BUF_202 (c2670_wire_354, G81_net_0);
bufg #(0, 0) BUF_203 (c2670_wire_340, G82_net_0);
bufg #(0, 0) BUF_204 (c2670_wire_313, G83_net_0);
notg #(0, 0) NOT_192 (c2670_wire_981, c2670_wire_435);
bufg #(0, 0) BUF_205 (c2670_wire_366, G84_net_0);
bufg #(0, 0) BUF_206 (c2670_wire_295, G85_net_0);
bufg #(0, 0) BUF_207 (c2670_wire_945, G86_net_0);
bufg #(0, 0) BUF_208 (c2670_wire_273, G87_net_0);
bufg #(0, 0) BUF_209 (c2670_wire_247, G88_net_0);
bufg #(0, 0) BUF_210 (c2670_wire_229, G89_net_0);
bufg #(0, 0) BUF_211 (c2670_wire_753, G9_net_0);
bufg #(0, 0) BUF_212 (c2670_wire_204, G90_net_0);
nor_n #(2, 0, 0) NOR_81 (c2670_wire_377, {c2670_wire_483_4, c2670_wire_489_6});
bufg #(0, 0) BUF_213 (c2670_wire_357, G91_net_0);
nor_n #(2, 0, 0) NOR_82 (c2670_wire_381, {c2670_wire_525_4, c2670_wire_552_6});
bufg #(0, 0) BUF_214 (c2670_wire_343, G92_net_0);
bufg #(0, 0) BUF_215 (c2670_wire_316, G93_net_0);
bufg #(0, 0) BUF_216 (c2670_wire_369, G94_net_0);
bufg #(0, 0) BUF_217 (c2670_wire_290, G95_net_0);
nor_n #(2, 0, 0) NOR_83 (c2670_wire_391, {c2670_wire_347_7, c2670_wire_574_5});
bufg #(0, 0) BUF_218 (c2670_wire_941, G96_net_0);
nor_n #(2, 0, 0) NOR_84 (c2670_wire_395, {c2670_wire_216_7, c2670_wire_234_7});
bufg #(0, 0) BUF_219 (c2670_wire_268, G97_net_0);
bufg #(0, 0) BUF_220 (c2670_wire_242, G98_net_0);
nor_n #(2, 0, 0) NOR_85 (c2670_wire_398, {c2670_wire_465_4, c2670_wire_466_4});
nor_n #(2, 0, 0) NOR_86 (c2670_wire_403, {c2670_wire_284_7, c2670_wire_302_8});
nor_n #(2, 0, 0) NOR_87 (c2670_wire_408, {c2670_wire_477_6, c2670_wire_557_6});
bufg #(0, 0) BUF_221 (c2670_wire_224, G99_net_0);
and_n #(2, 0, 0) AND_330 (c2670_wire_420, {c2670_wire_981, c2670_wire_972});
or_n #(2, 0, 0) OR_191 (c2670_wire_431, {c2670_wire_442, c2670_wire_974});
and_n #(2, 0, 0) AND_331 (c2670_wire_568, {c2670_wire_429, c2670_wire_982});
or_n #(2, 0, 0) OR_192 (c2670_wire_982, {c2670_wire_445, c2670_wire_976});

endmodule
