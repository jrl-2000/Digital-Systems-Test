/****************************************************************************
 *                                                                          *
 *  FLAT VERSION of HIGH-LEVEL MODEL for c2670                              *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *  Verified  by: Jonathan David Hauke (jhauke@eecs.umich.edu)              *
 *                                                                          *
 *                Oct 20, 1998                                              *
 *                                                                          *
****************************************************************************/
// Flat Verilog File 
module c2670g (
	in81, in92, in91, in90, in89, in88, in87, 
	in86, in85, in93, in43, in54, in53, in52, in51, 
	in50, in49, in48, in47, in55, in56, in66, in65, 
	in64, in63, in62, in61, in60, in67, in68, in79, 
	in78, in77, in76, in75, in74, in73, in72, in80, 
	in131, in141, in140, in139, in138, in137, in136, in135, 
	in142, in95, in105, in104, in103, in102, in101, in100, 
	in99, in106, in119, in129, in128, in127, in126, in125, 
	in124, in123, in130, in107, in117, in116, in115, in114, 
	in113, in112, in111, in118, in1971, in1966, in1961, in1956, 
	in1348, in1341, in2090, in2084, in2078, in2072, in2067, in1996, 
	in1991, in1986, in1981, in1976, in2096, in2100, in2678, in2474, 
	in2427, in2430, in2451, in2454, in2443, in2446, in2435, in2438, 
	in24, in6, in23, in22, in21, in5, in20, in4, 
	in19, in28, in35, in34, in27, in33, in26, in32, 
	in25, in651, in543, in2105, in2104, in1384, in40, in16, 
	in29, in11, in8, in37, in14, in44, in132, in82, 
	in96, in69, in120, in57, in108, in2106, in567, in559, 
	in860, in868, in452, in2066, in1083, in94, in7, in661, 
	in1, in2, in3, in15, in36, in483, in169, in174, 
	in177, in178, in179, in180, in181, in182, in183, in184, 
	in185, in186, in189, in190, in191, in192, in193, in194, 
	in195, in196, in197, in198, in199, in200, in201, in202, 
	in203, in204, in205, in206, in207, in208, in209, in210, 
	in211, in212, in213, in214, in215, in239, in240, in241, 
	in242, in243, in244, in245, in246, in247, in248, in249, 
	in250, in251, in252, in253, in254, in255, in256, in257, 
	in262, in263, in264, in265, in266, in267, in268, in269, 
	in270, in271, in272, in273, in274, in275, in276, in277, 
	in278, in279,
	out329, out231, out311, out150, out308, out225, out395, 
	out397, out227, out229, out401, out319, out325, out261, out220, 
	out221, out219, out218, out235, out236, out237, out238, out335, 
	out350, out391, out409, out337, out384, out411, out367, out369, 
	out173, out295, out331, out145, out148, out282, out323, out284, 
	out321, out297, out280, out153, out290, out305, out288, out303, 
	out286, out301, out299, out166, out168, out171, out162, out160, 
	out164, out156, out223, out217, out234, out259, out176, out188, 
	out158, out169, out174, out177, out178, out179, out180, out181, 
	out182, out183, out184, out185, out186, out189, out190, out191, 
	out192, out193, out194, out195, out196, out197, out198, out199, 
	out200, out201, out202, out203, out204, out205, out206, out207, 
	out208, out209, out210, out211, out212, out213, out214, out215, 
	out239, out240, out241, out242, out243, out244, out245, out246, 
	out247, out248, out249, out250, out251, out252, out253, out254, 
	out255, out256, out257, out262, out263, out264, out265, out266, 
	out267, out268, out269, out270, out271, out272, out273, out274, 
	out275, out276, out277, out278, out279);

   input
	in81, in92, in91, in90, in89, in88, in87, 
	in86, in85, in93, in43, in54, in53, in52, in51, 
	in50, in49, in48, in47, in55, in56, in66, in65, 
	in64, in63, in62, in61, in60, in67, in68, in79, 
	in78, in77, in76, in75, in74, in73, in72, in80, 
	in131, in141, in140, in139, in138, in137, in136, in135, 
	in142, in95, in105, in104, in103, in102, in101, in100, 
	in99, in106, in119, in129, in128, in127, in126, in125, 
	in124, in123, in130, in107, in117, in116, in115, in114, 
	in113, in112, in111, in118, in1971, in1966, in1961, in1956, 
	in1348, in1341, in2090, in2084, in2078, in2072, in2067, in1996, 
	in1991, in1986, in1981, in1976, in2096, in2100, in2678, in2474, 
	in2427, in2430, in2451, in2454, in2443, in2446, in2435, in2438, 
	in24, in6, in23, in22, in21, in5, in20, in4, 
	in19, in28, in35, in34, in27, in33, in26, in32, 
	in25, in651, in543, in2105, in2104, in1384, in40, in16, 
	in29, in11, in8, in37, in14, in44, in132, in82, 
	in96, in69, in120, in57, in108, in2106, in567, in559, 
	in860, in868, in452, in2066, in1083, in94, in7, in661, 
	in1, in2, in3, in15, in36, in483, in169, in174, 
	in177, in178, in179, in180, in181, in182, in183, in184, 
	in185, in186, in189, in190, in191, in192, in193, in194, 
	in195, in196, in197, in198, in199, in200, in201, in202, 
	in203, in204, in205, in206, in207, in208, in209, in210, 
	in211, in212, in213, in214, in215, in239, in240, in241, 
	in242, in243, in244, in245, in246, in247, in248, in249, 
	in250, in251, in252, in253, in254, in255, in256, in257, 
	in262, in263, in264, in265, in266, in267, in268, in269, 
	in270, in271, in272, in273, in274, in275, in276, in277, 
	in278, in279;

   output
	out329, out231, out311, out150, out308, out225, out395, 
	out397, out227, out229, out401, out319, out325, out261, out220, 
	out221, out219, out218, out235, out236, out237, out238, out335, 
	out350, out391, out409, out337, out384, out411, out367, out369, 
	out173, out295, out331, out145, out148, out282, out323, out284, 
	out321, out297, out280, out153, out290, out305, out288, out303, 
	out286, out301, out299, out166, out168, out171, out162, out160, 
	out164, out156, out223, out217, out234, out259, out176, out188, 
	out158, out169, out174, out177, out178, out179, out180, out181, 
	out182, out183, out184, out185, out186, out189, out190, out191, 
	out192, out193, out194, out195, out196, out197, out198, out199, 
	out200, out201, out202, out203, out204, out205, out206, out207, 
	out208, out209, out210, out211, out212, out213, out214, out215, 
	out239, out240, out241, out242, out243, out244, out245, out246, 
	out247, out248, out249, out250, out251, out252, out253, out254, 
	out255, out256, out257, out262, out263, out264, out265, out266, 
	out267, out268, out269, out270, out271, out272, out273, out274, 
	out275, out276, out277, out278, out279;

inv M1_Mux0_Mux0(in651, M1_Mux0_Not_Cont0);
inv M1_Mux0_Mux1(in543, M1_Mux0_Not_Cont1);
and3 M1_Mux0_Mux2(in81, M1_Mux0_Not_Cont0, M1_Mux0_Not_Cont1, M1_Mux0_line2);
and3 M1_Mux0_Mux3(in43, M1_Mux0_Not_Cont0, in543, M1_Mux0_line3);
and3 M1_Mux0_Mux4(in56, in651, M1_Mux0_Not_Cont1, M1_Mux0_line4);
and3 M1_Mux0_Mux5(in68, in651, in543, M1_Mux0_line5);
or4 M1_Mux0_Mux6(M1_Mux0_line2, M1_Mux0_line3, M1_Mux0_line4, M1_Mux0_line5, Abus_0);
inv M1_Mux1_Mux0(in651, M1_Mux1_Not_Cont0);
inv M1_Mux1_Mux1(in543, M1_Mux1_Not_Cont1);
and3 M1_Mux1_Mux2(in92, M1_Mux1_Not_Cont0, M1_Mux1_Not_Cont1, M1_Mux1_line2);
and3 M1_Mux1_Mux3(in54, M1_Mux1_Not_Cont0, in543, M1_Mux1_line3);
and3 M1_Mux1_Mux4(in66, in651, M1_Mux1_Not_Cont1, M1_Mux1_line4);
and3 M1_Mux1_Mux5(in79, in651, in543, M1_Mux1_line5);
or4 M1_Mux1_Mux6(M1_Mux1_line2, M1_Mux1_line3, M1_Mux1_line4, M1_Mux1_line5, Abus_1);
inv M1_Mux2_Mux0(in651, M1_Mux2_Not_Cont0);
inv M1_Mux2_Mux1(in543, M1_Mux2_Not_Cont1);
and3 M1_Mux2_Mux2(in91, M1_Mux2_Not_Cont0, M1_Mux2_Not_Cont1, M1_Mux2_line2);
and3 M1_Mux2_Mux3(in53, M1_Mux2_Not_Cont0, in543, M1_Mux2_line3);
and3 M1_Mux2_Mux4(in65, in651, M1_Mux2_Not_Cont1, M1_Mux2_line4);
and3 M1_Mux2_Mux5(in78, in651, in543, M1_Mux2_line5);
or4 M1_Mux2_Mux6(M1_Mux2_line2, M1_Mux2_line3, M1_Mux2_line4, M1_Mux2_line5, Abus_2);
inv M1_Mux3_Mux0(in651, M1_Mux3_Not_Cont0);
inv M1_Mux3_Mux1(in543, M1_Mux3_Not_Cont1);
and3 M1_Mux3_Mux2(in90, M1_Mux3_Not_Cont0, M1_Mux3_Not_Cont1, M1_Mux3_line2);
and3 M1_Mux3_Mux3(in52, M1_Mux3_Not_Cont0, in543, M1_Mux3_line3);
and3 M1_Mux3_Mux4(in64, in651, M1_Mux3_Not_Cont1, M1_Mux3_line4);
and3 M1_Mux3_Mux5(in77, in651, in543, M1_Mux3_line5);
or4 M1_Mux3_Mux6(M1_Mux3_line2, M1_Mux3_line3, M1_Mux3_line4, M1_Mux3_line5, Abus_3);
inv M1_Mux4_Mux0(in651, M1_Mux4_Not_Cont0);
inv M1_Mux4_Mux1(in543, M1_Mux4_Not_Cont1);
and3 M1_Mux4_Mux2(in89, M1_Mux4_Not_Cont0, M1_Mux4_Not_Cont1, M1_Mux4_line2);
and3 M1_Mux4_Mux3(in51, M1_Mux4_Not_Cont0, in543, M1_Mux4_line3);
and3 M1_Mux4_Mux4(in63, in651, M1_Mux4_Not_Cont1, M1_Mux4_line4);
and3 M1_Mux4_Mux5(in76, in651, in543, M1_Mux4_line5);
or4 M1_Mux4_Mux6(M1_Mux4_line2, M1_Mux4_line3, M1_Mux4_line4, M1_Mux4_line5, Abus_4);
inv M1_Mux5_Mux0(in651, M1_Mux5_Not_Cont0);
inv M1_Mux5_Mux1(in543, M1_Mux5_Not_Cont1);
and3 M1_Mux5_Mux2(in88, M1_Mux5_Not_Cont0, M1_Mux5_Not_Cont1, M1_Mux5_line2);
and3 M1_Mux5_Mux3(in50, M1_Mux5_Not_Cont0, in543, M1_Mux5_line3);
and3 M1_Mux5_Mux4(in62, in651, M1_Mux5_Not_Cont1, M1_Mux5_line4);
and3 M1_Mux5_Mux5(in75, in651, in543, M1_Mux5_line5);
or4 M1_Mux5_Mux6(M1_Mux5_line2, M1_Mux5_line3, M1_Mux5_line4, M1_Mux5_line5, Abus_5);
inv M1_Mux6_Mux0(in651, M1_Mux6_Not_Cont0);
inv M1_Mux6_Mux1(in543, M1_Mux6_Not_Cont1);
and3 M1_Mux6_Mux2(in87, M1_Mux6_Not_Cont0, M1_Mux6_Not_Cont1, M1_Mux6_line2);
and3 M1_Mux6_Mux3(in49, M1_Mux6_Not_Cont0, in543, M1_Mux6_line3);
and3 M1_Mux6_Mux4(vdd, in651, M1_Mux6_Not_Cont1, M1_Mux6_line4);
and3 M1_Mux6_Mux5(in74, in651, in543, M1_Mux6_line5);
or4 M1_Mux6_Mux6(M1_Mux6_line2, M1_Mux6_line3, M1_Mux6_line4, M1_Mux6_line5, Abus_6);
inv M1_Mux7_Mux0(in651, M1_Mux7_Not_Cont0);
inv M1_Mux7_Mux1(in543, M1_Mux7_Not_Cont1);
and3 M1_Mux7_Mux2(in86, M1_Mux7_Not_Cont0, M1_Mux7_Not_Cont1, M1_Mux7_line2);
and3 M1_Mux7_Mux3(in48, M1_Mux7_Not_Cont0, in543, M1_Mux7_line3);
and3 M1_Mux7_Mux4(in61, in651, M1_Mux7_Not_Cont1, M1_Mux7_line4);
and3 M1_Mux7_Mux5(in73, in651, in543, M1_Mux7_line5);
or4 M1_Mux7_Mux6(M1_Mux7_line2, M1_Mux7_line3, M1_Mux7_line4, M1_Mux7_line5, Abus_7);
inv M1_Mux8_Mux0(in651, M1_Mux8_Not_Cont0);
inv M1_Mux8_Mux1(in543, M1_Mux8_Not_Cont1);
and3 M1_Mux8_Mux2(in85, M1_Mux8_Not_Cont0, M1_Mux8_Not_Cont1, M1_Mux8_line2);
and3 M1_Mux8_Mux3(in47, M1_Mux8_Not_Cont0, in543, M1_Mux8_line3);
and3 M1_Mux8_Mux4(in60, in651, M1_Mux8_Not_Cont1, M1_Mux8_line4);
and3 M1_Mux8_Mux5(in72, in651, in543, M1_Mux8_line5);
or4 M1_Mux8_Mux6(M1_Mux8_line2, M1_Mux8_line3, M1_Mux8_line4, M1_Mux8_line5, Abus_8);
inv M1_Mux9_Mux0(in651, M1_Mux9_Not_Cont0);
inv M1_Mux9_Mux1(in543, M1_Mux9_Not_Cont1);
and3 M1_Mux9_Mux2(in93, M1_Mux9_Not_Cont0, M1_Mux9_Not_Cont1, M1_Mux9_line2);
and3 M1_Mux9_Mux3(in55, M1_Mux9_Not_Cont0, in543, M1_Mux9_line3);
and3 M1_Mux9_Mux4(in67, in651, M1_Mux9_Not_Cont1, M1_Mux9_line4);
and3 M1_Mux9_Mux5(in80, in651, in543, M1_Mux9_line5);
or4 M1_Mux9_Mux6(M1_Mux9_line2, M1_Mux9_line3, M1_Mux9_line4, M1_Mux9_line5, Abus_9);
inv M2_Mux0_Mux0(in2105, M2_Mux0_Not_Cont0);
inv M2_Mux0_Mux1(in2104, M2_Mux0_Not_Cont1);
and3 M2_Mux0_Mux2(in131, M2_Mux0_Not_Cont0, M2_Mux0_Not_Cont1, M2_Mux0_line2);
and3 M2_Mux0_Mux3(in95, M2_Mux0_Not_Cont0, in2104, M2_Mux0_line3);
and3 M2_Mux0_Mux4(in119, in2105, M2_Mux0_Not_Cont1, M2_Mux0_line4);
and3 M2_Mux0_Mux5(in107, in2105, in2104, M2_Mux0_line5);
or4 M2_Mux0_Mux6(M2_Mux0_line2, M2_Mux0_line3, M2_Mux0_line4, M2_Mux0_line5, Bbus_0);
inv M2_Mux1_Mux0(in2105, M2_Mux1_Not_Cont0);
inv M2_Mux1_Mux1(in2104, M2_Mux1_Not_Cont1);
and3 M2_Mux1_Mux2(in141, M2_Mux1_Not_Cont0, M2_Mux1_Not_Cont1, M2_Mux1_line2);
and3 M2_Mux1_Mux3(in105, M2_Mux1_Not_Cont0, in2104, M2_Mux1_line3);
and3 M2_Mux1_Mux4(in129, in2105, M2_Mux1_Not_Cont1, M2_Mux1_line4);
and3 M2_Mux1_Mux5(in117, in2105, in2104, M2_Mux1_line5);
or4 M2_Mux1_Mux6(M2_Mux1_line2, M2_Mux1_line3, M2_Mux1_line4, M2_Mux1_line5, Bbus_1);
inv M2_Mux2_Mux0(in2105, M2_Mux2_Not_Cont0);
inv M2_Mux2_Mux1(in2104, M2_Mux2_Not_Cont1);
and3 M2_Mux2_Mux2(in140, M2_Mux2_Not_Cont0, M2_Mux2_Not_Cont1, M2_Mux2_line2);
and3 M2_Mux2_Mux3(in104, M2_Mux2_Not_Cont0, in2104, M2_Mux2_line3);
and3 M2_Mux2_Mux4(in128, in2105, M2_Mux2_Not_Cont1, M2_Mux2_line4);
and3 M2_Mux2_Mux5(in116, in2105, in2104, M2_Mux2_line5);
or4 M2_Mux2_Mux6(M2_Mux2_line2, M2_Mux2_line3, M2_Mux2_line4, M2_Mux2_line5, Bbus_2);
inv M2_Mux3_Mux0(in2105, M2_Mux3_Not_Cont0);
inv M2_Mux3_Mux1(in2104, M2_Mux3_Not_Cont1);
and3 M2_Mux3_Mux2(in139, M2_Mux3_Not_Cont0, M2_Mux3_Not_Cont1, M2_Mux3_line2);
and3 M2_Mux3_Mux3(in103, M2_Mux3_Not_Cont0, in2104, M2_Mux3_line3);
and3 M2_Mux3_Mux4(in127, in2105, M2_Mux3_Not_Cont1, M2_Mux3_line4);
and3 M2_Mux3_Mux5(in115, in2105, in2104, M2_Mux3_line5);
or4 M2_Mux3_Mux6(M2_Mux3_line2, M2_Mux3_line3, M2_Mux3_line4, M2_Mux3_line5, Bbus_3);
inv M2_Mux4_Mux0(in2105, M2_Mux4_Not_Cont0);
inv M2_Mux4_Mux1(in2104, M2_Mux4_Not_Cont1);
and3 M2_Mux4_Mux2(in138, M2_Mux4_Not_Cont0, M2_Mux4_Not_Cont1, M2_Mux4_line2);
and3 M2_Mux4_Mux3(in102, M2_Mux4_Not_Cont0, in2104, M2_Mux4_line3);
and3 M2_Mux4_Mux4(in126, in2105, M2_Mux4_Not_Cont1, M2_Mux4_line4);
and3 M2_Mux4_Mux5(in114, in2105, in2104, M2_Mux4_line5);
or4 M2_Mux4_Mux6(M2_Mux4_line2, M2_Mux4_line3, M2_Mux4_line4, M2_Mux4_line5, Bbus_4);
inv M2_Mux5_Mux0(in2105, M2_Mux5_Not_Cont0);
inv M2_Mux5_Mux1(in2104, M2_Mux5_Not_Cont1);
and3 M2_Mux5_Mux2(in137, M2_Mux5_Not_Cont0, M2_Mux5_Not_Cont1, M2_Mux5_line2);
and3 M2_Mux5_Mux3(in101, M2_Mux5_Not_Cont0, in2104, M2_Mux5_line3);
and3 M2_Mux5_Mux4(in125, in2105, M2_Mux5_Not_Cont1, M2_Mux5_line4);
and3 M2_Mux5_Mux5(in113, in2105, in2104, M2_Mux5_line5);
or4 M2_Mux5_Mux6(M2_Mux5_line2, M2_Mux5_line3, M2_Mux5_line4, M2_Mux5_line5, Bbus_5);
inv M2_Mux6_Mux0(in2105, M2_Mux6_Not_Cont0);
inv M2_Mux6_Mux1(in2104, M2_Mux6_Not_Cont1);
and3 M2_Mux6_Mux2(in136, M2_Mux6_Not_Cont0, M2_Mux6_Not_Cont1, M2_Mux6_line2);
and3 M2_Mux6_Mux3(in100, M2_Mux6_Not_Cont0, in2104, M2_Mux6_line3);
and3 M2_Mux6_Mux4(in124, in2105, M2_Mux6_Not_Cont1, M2_Mux6_line4);
and3 M2_Mux6_Mux5(in112, in2105, in2104, M2_Mux6_line5);
or4 M2_Mux6_Mux6(M2_Mux6_line2, M2_Mux6_line3, M2_Mux6_line4, M2_Mux6_line5, Bbus_6);
inv M2_Mux7_Mux0(in2105, M2_Mux7_Not_Cont0);
inv M2_Mux7_Mux1(in2104, M2_Mux7_Not_Cont1);
and3 M2_Mux7_Mux2(in135, M2_Mux7_Not_Cont0, M2_Mux7_Not_Cont1, M2_Mux7_line2);
and3 M2_Mux7_Mux3(in99, M2_Mux7_Not_Cont0, in2104, M2_Mux7_line3);
and3 M2_Mux7_Mux4(in123, in2105, M2_Mux7_Not_Cont1, M2_Mux7_line4);
and3 M2_Mux7_Mux5(in111, in2105, in2104, M2_Mux7_line5);
or4 M2_Mux7_Mux6(M2_Mux7_line2, M2_Mux7_line3, M2_Mux7_line4, M2_Mux7_line5, Bbus_7);
inv M2_Mux8_Mux0(in2105, M2_Mux8_Not_Cont0);
inv M2_Mux8_Mux1(in2104, M2_Mux8_Not_Cont1);
and3 M2_Mux8_Mux2(in142, M2_Mux8_Not_Cont0, M2_Mux8_Not_Cont1, M2_Mux8_line2);
and3 M2_Mux8_Mux3(in106, M2_Mux8_Not_Cont0, in2104, M2_Mux8_line3);
and3 M2_Mux8_Mux4(in130, in2105, M2_Mux8_Not_Cont1, M2_Mux8_line4);
and3 M2_Mux8_Mux5(in118, in2105, in2104, M2_Mux8_line5);
or4 M2_Mux8_Mux6(M2_Mux8_line2, M2_Mux8_line3, M2_Mux8_line4, M2_Mux8_line5, Bbus_8);
inv M2_Mux9_Mux0(in2105, M2_Mux9_Not_Cont0);
inv M2_Mux9_Mux1(in2104, M2_Mux9_Not_Cont1);
and3 M2_Mux9_Mux2(vdd, M2_Mux9_Not_Cont0, M2_Mux9_Not_Cont1, M2_Mux9_line2);
and3 M2_Mux9_Mux3(vdd, M2_Mux9_Not_Cont0, in2104, M2_Mux9_line3);
and3 M2_Mux9_Mux4(vdd, in2105, M2_Mux9_Not_Cont1, M2_Mux9_line4);
and3 M2_Mux9_Mux5(vdd, in2105, in2104, M2_Mux9_line5);
or4 M2_Mux9_Mux6(M2_Mux9_line2, M2_Mux9_line3, M2_Mux9_line4, M2_Mux9_line5, Bbus_9);
inv M3_UM3_0(Bbus_5, M3_NotB5);
inv M3_UM3_1(in1384, M3_NotMask1);
and2 M3_UM3_2(Bbus_4, M3_NotMask1, M3_line2);
and3 M3_UM3_3(M3_NotB5, M3_line2, in40, ContAlpha);
inv M3_UM3_4(M3_line2, M3_line4);
and3 M3_UM3_5(in40, M3_line4, M3_NotB5, ContBeta);
and2 M4_UM4_0_MB0(Abus_4, in8, M4_XMbus_4);
and2 M4_UM4_0_MB1(Abus_5, in8, M4_XMbus_5);
inv M4_UM4_0_MB2(ContAlpha, M4_UM4_0_NotAlpha);
and2 M4_UM4_0_MB3(Abus_6, M4_UM4_0_NotAlpha, M4_UM4_0_line3);
and2 M4_UM4_0_MB4(M4_UM4_0_line3, in8, M4_XMbus_6);
and2 M4_UM4_0_MB5(Abus_7, M4_UM4_0_NotAlpha, M4_UM4_0_line5);
and2 M4_UM4_0_MB6(M4_UM4_0_line5, in8, M4_XMbus_7);
and2 M4_UM4_0_MB7(Abus_8, M4_UM4_0_NotAlpha, M4_UM4_0_line7);
and2 M4_UM4_0_MB8(M4_UM4_0_line7, ContBeta, M4_XMbus_8);
and2 M4_UM4_0_MB9(Bbus_0, M4_UM4_0_NotAlpha, M4_UM4_0_line9);
and2 M4_UM4_0_MB10(M4_UM4_0_line9, ContBeta, M4_XMbus_9);
and2 M4_UM4_0_MB11(Bbus_1, M4_UM4_0_NotAlpha, M4_UM4_0_line11);
and2 M4_UM4_0_MB12(M4_UM4_0_line11, ContBeta, M4_XMbus_10);
and2 M4_UM4_0_MB13(Bbus_2, M4_UM4_0_NotAlpha, M4_UM4_0_line13);
and2 M4_UM4_0_MB14(M4_UM4_0_line13, ContBeta, M4_XMbus_11);
and2 M4_UM4_1_MB0(Ybus_4, in8, M4_YMbus_4);
and2 M4_UM4_1_MB1(Ybus_5, in8, M4_YMbus_5);
inv M4_UM4_1_MB2(ContAlpha, M4_UM4_1_NotAlpha);
and2 M4_UM4_1_MB3(Ybus_6, M4_UM4_1_NotAlpha, M4_UM4_1_line3);
and2 M4_UM4_1_MB4(M4_UM4_1_line3, in8, M4_YMbus_6);
and2 M4_UM4_1_MB5(Ybus_7, M4_UM4_1_NotAlpha, M4_UM4_1_line5);
and2 M4_UM4_1_MB6(M4_UM4_1_line5, in8, M4_YMbus_7);
and2 M4_UM4_1_MB7(Ybus_8, M4_UM4_1_NotAlpha, M4_UM4_1_line7);
and2 M4_UM4_1_MB8(M4_UM4_1_line7, ContBeta, M4_YMbus_8);
and2 M4_UM4_1_MB9(Ybus_9, M4_UM4_1_NotAlpha, M4_UM4_1_line9);
and2 M4_UM4_1_MB10(M4_UM4_1_line9, ContBeta, M4_YMbus_9);
and2 M4_UM4_1_MB11(Ybus_10, M4_UM4_1_NotAlpha, M4_UM4_1_line11);
and2 M4_UM4_1_MB12(M4_UM4_1_line11, ContBeta, M4_YMbus_10);
and2 M4_UM4_1_MB13(Ybus_11, M4_UM4_1_NotAlpha, M4_UM4_1_line13);
and2 M4_UM4_1_MB14(M4_UM4_1_line13, ContBeta, M4_YMbus_11);
inv M4_UM4_2_Inv12_0(Abus_0, M4_Not_XMbus_0);
inv M4_UM4_2_Inv12_1(Abus_1, M4_Not_XMbus_1);
inv M4_UM4_2_Inv12_2(Abus_2, M4_Not_XMbus_2);
inv M4_UM4_2_Inv12_3(Abus_3, M4_Not_XMbus_3);
inv M4_UM4_2_Inv12_4(M4_XMbus_4, M4_Not_XMbus_4);
inv M4_UM4_2_Inv12_5(M4_XMbus_5, M4_Not_XMbus_5);
inv M4_UM4_2_Inv12_6(M4_XMbus_6, M4_Not_XMbus_6);
inv M4_UM4_2_Inv12_7(M4_XMbus_7, M4_Not_XMbus_7);
inv M4_UM4_2_Inv12_8(M4_XMbus_8, M4_Not_XMbus_8);
inv M4_UM4_2_Inv12_9(M4_XMbus_9, M4_Not_XMbus_9);
inv M4_UM4_2_Inv12_10(M4_XMbus_10, M4_Not_XMbus_10);
inv M4_UM4_2_Inv12_11(M4_XMbus_11, M4_Not_XMbus_11);
and2 M4_UM4_3_GP_CalGP0(M4_Not_XMbus_0, Ybus_0, M4_UM4_3_Gbus_0);
and2 M4_UM4_3_GP_CalGP1(M4_Not_XMbus_1, Ybus_1, M4_UM4_3_Gbus_1);
and2 M4_UM4_3_GP_CalGP2(M4_Not_XMbus_2, Ybus_2, M4_UM4_3_Gbus_2);
and2 M4_UM4_3_GP_CalGP3(M4_Not_XMbus_3, Ybus_3, M4_UM4_3_Gbus_3);
and2 M4_UM4_3_GP_CalGP4(M4_Not_XMbus_4, M4_YMbus_4, M4_UM4_3_Gbus_4);
and2 M4_UM4_3_GP_CalGP5(M4_Not_XMbus_5, M4_YMbus_5, M4_UM4_3_Gbus_5);
and2 M4_UM4_3_GP_CalGP6(M4_Not_XMbus_6, M4_YMbus_6, M4_UM4_3_Gbus_6);
and2 M4_UM4_3_GP_CalGP7(M4_Not_XMbus_7, M4_YMbus_7, M4_UM4_3_Gbus_7);
and2 M4_UM4_3_GP_CalGP8(M4_Not_XMbus_8, M4_YMbus_8, M4_UM4_3_Gbus_8);
and2 M4_UM4_3_GP_CalGP9(M4_Not_XMbus_9, M4_YMbus_9, M4_UM4_3_Gbus_9);
and2 M4_UM4_3_GP_CalGP10(M4_Not_XMbus_10, M4_YMbus_10, M4_UM4_3_Gbus_10);
and2 M4_UM4_3_GP_CalGP11(M4_Not_XMbus_11, M4_YMbus_11, M4_UM4_3_Gbus_11);
inv M4_UM4_3_GP_CalGP12_Xo0(M4_Not_XMbus_0, M4_UM4_3_GP_CalGP12_NotA);
inv M4_UM4_3_GP_CalGP12_Xo1(Ybus_0, M4_UM4_3_GP_CalGP12_NotB);
nand2 M4_UM4_3_GP_CalGP12_Xo2(M4_UM4_3_GP_CalGP12_NotA, Ybus_0, M4_UM4_3_GP_CalGP12_line2);
nand2 M4_UM4_3_GP_CalGP12_Xo3(M4_UM4_3_GP_CalGP12_NotB, M4_Not_XMbus_0, M4_UM4_3_GP_CalGP12_line3);
nand2 M4_UM4_3_GP_CalGP12_Xo4(M4_UM4_3_GP_CalGP12_line2, M4_UM4_3_GP_CalGP12_line3, M4_UM4_3_Pbus_0);
inv M4_UM4_3_GP_CalGP13_Xo0(M4_Not_XMbus_1, M4_UM4_3_GP_CalGP13_NotA);
inv M4_UM4_3_GP_CalGP13_Xo1(Ybus_1, M4_UM4_3_GP_CalGP13_NotB);
nand2 M4_UM4_3_GP_CalGP13_Xo2(M4_UM4_3_GP_CalGP13_NotA, Ybus_1, M4_UM4_3_GP_CalGP13_line2);
nand2 M4_UM4_3_GP_CalGP13_Xo3(M4_UM4_3_GP_CalGP13_NotB, M4_Not_XMbus_1, M4_UM4_3_GP_CalGP13_line3);
nand2 M4_UM4_3_GP_CalGP13_Xo4(M4_UM4_3_GP_CalGP13_line2, M4_UM4_3_GP_CalGP13_line3, M4_UM4_3_Pbus_1);
inv M4_UM4_3_GP_CalGP14_Xo0(M4_Not_XMbus_2, M4_UM4_3_GP_CalGP14_NotA);
inv M4_UM4_3_GP_CalGP14_Xo1(Ybus_2, M4_UM4_3_GP_CalGP14_NotB);
nand2 M4_UM4_3_GP_CalGP14_Xo2(M4_UM4_3_GP_CalGP14_NotA, Ybus_2, M4_UM4_3_GP_CalGP14_line2);
nand2 M4_UM4_3_GP_CalGP14_Xo3(M4_UM4_3_GP_CalGP14_NotB, M4_Not_XMbus_2, M4_UM4_3_GP_CalGP14_line3);
nand2 M4_UM4_3_GP_CalGP14_Xo4(M4_UM4_3_GP_CalGP14_line2, M4_UM4_3_GP_CalGP14_line3, M4_UM4_3_Pbus_2);
inv M4_UM4_3_GP_CalGP15_Xo0(M4_Not_XMbus_3, M4_UM4_3_GP_CalGP15_NotA);
inv M4_UM4_3_GP_CalGP15_Xo1(Ybus_3, M4_UM4_3_GP_CalGP15_NotB);
nand2 M4_UM4_3_GP_CalGP15_Xo2(M4_UM4_3_GP_CalGP15_NotA, Ybus_3, M4_UM4_3_GP_CalGP15_line2);
nand2 M4_UM4_3_GP_CalGP15_Xo3(M4_UM4_3_GP_CalGP15_NotB, M4_Not_XMbus_3, M4_UM4_3_GP_CalGP15_line3);
nand2 M4_UM4_3_GP_CalGP15_Xo4(M4_UM4_3_GP_CalGP15_line2, M4_UM4_3_GP_CalGP15_line3, M4_UM4_3_Pbus_3);
inv M4_UM4_3_GP_CalGP16_Xo0(M4_Not_XMbus_4, M4_UM4_3_GP_CalGP16_NotA);
inv M4_UM4_3_GP_CalGP16_Xo1(M4_YMbus_4, M4_UM4_3_GP_CalGP16_NotB);
nand2 M4_UM4_3_GP_CalGP16_Xo2(M4_UM4_3_GP_CalGP16_NotA, M4_YMbus_4, M4_UM4_3_GP_CalGP16_line2);
nand2 M4_UM4_3_GP_CalGP16_Xo3(M4_UM4_3_GP_CalGP16_NotB, M4_Not_XMbus_4, M4_UM4_3_GP_CalGP16_line3);
nand2 M4_UM4_3_GP_CalGP16_Xo4(M4_UM4_3_GP_CalGP16_line2, M4_UM4_3_GP_CalGP16_line3, M4_UM4_3_Pbus_4);
inv M4_UM4_3_GP_CalGP17_Xo0(M4_Not_XMbus_5, M4_UM4_3_GP_CalGP17_NotA);
inv M4_UM4_3_GP_CalGP17_Xo1(M4_YMbus_5, M4_UM4_3_GP_CalGP17_NotB);
nand2 M4_UM4_3_GP_CalGP17_Xo2(M4_UM4_3_GP_CalGP17_NotA, M4_YMbus_5, M4_UM4_3_GP_CalGP17_line2);
nand2 M4_UM4_3_GP_CalGP17_Xo3(M4_UM4_3_GP_CalGP17_NotB, M4_Not_XMbus_5, M4_UM4_3_GP_CalGP17_line3);
nand2 M4_UM4_3_GP_CalGP17_Xo4(M4_UM4_3_GP_CalGP17_line2, M4_UM4_3_GP_CalGP17_line3, M4_UM4_3_Pbus_5);
inv M4_UM4_3_GP_CalGP18_Xo0(M4_Not_XMbus_6, M4_UM4_3_GP_CalGP18_NotA);
inv M4_UM4_3_GP_CalGP18_Xo1(M4_YMbus_6, M4_UM4_3_GP_CalGP18_NotB);
nand2 M4_UM4_3_GP_CalGP18_Xo2(M4_UM4_3_GP_CalGP18_NotA, M4_YMbus_6, M4_UM4_3_GP_CalGP18_line2);
nand2 M4_UM4_3_GP_CalGP18_Xo3(M4_UM4_3_GP_CalGP18_NotB, M4_Not_XMbus_6, M4_UM4_3_GP_CalGP18_line3);
nand2 M4_UM4_3_GP_CalGP18_Xo4(M4_UM4_3_GP_CalGP18_line2, M4_UM4_3_GP_CalGP18_line3, M4_UM4_3_Pbus_6);
inv M4_UM4_3_GP_CalGP19_Xo0(M4_Not_XMbus_7, M4_UM4_3_GP_CalGP19_NotA);
inv M4_UM4_3_GP_CalGP19_Xo1(M4_YMbus_7, M4_UM4_3_GP_CalGP19_NotB);
nand2 M4_UM4_3_GP_CalGP19_Xo2(M4_UM4_3_GP_CalGP19_NotA, M4_YMbus_7, M4_UM4_3_GP_CalGP19_line2);
nand2 M4_UM4_3_GP_CalGP19_Xo3(M4_UM4_3_GP_CalGP19_NotB, M4_Not_XMbus_7, M4_UM4_3_GP_CalGP19_line3);
nand2 M4_UM4_3_GP_CalGP19_Xo4(M4_UM4_3_GP_CalGP19_line2, M4_UM4_3_GP_CalGP19_line3, M4_UM4_3_Pbus_7);
inv M4_UM4_3_GP_CalGP20_Xo0(M4_Not_XMbus_8, M4_UM4_3_GP_CalGP20_NotA);
inv M4_UM4_3_GP_CalGP20_Xo1(M4_YMbus_8, M4_UM4_3_GP_CalGP20_NotB);
nand2 M4_UM4_3_GP_CalGP20_Xo2(M4_UM4_3_GP_CalGP20_NotA, M4_YMbus_8, M4_UM4_3_GP_CalGP20_line2);
nand2 M4_UM4_3_GP_CalGP20_Xo3(M4_UM4_3_GP_CalGP20_NotB, M4_Not_XMbus_8, M4_UM4_3_GP_CalGP20_line3);
nand2 M4_UM4_3_GP_CalGP20_Xo4(M4_UM4_3_GP_CalGP20_line2, M4_UM4_3_GP_CalGP20_line3, M4_UM4_3_Pbus_8);
inv M4_UM4_3_GP_CalGP21_Xo0(M4_Not_XMbus_9, M4_UM4_3_GP_CalGP21_NotA);
inv M4_UM4_3_GP_CalGP21_Xo1(M4_YMbus_9, M4_UM4_3_GP_CalGP21_NotB);
nand2 M4_UM4_3_GP_CalGP21_Xo2(M4_UM4_3_GP_CalGP21_NotA, M4_YMbus_9, M4_UM4_3_GP_CalGP21_line2);
nand2 M4_UM4_3_GP_CalGP21_Xo3(M4_UM4_3_GP_CalGP21_NotB, M4_Not_XMbus_9, M4_UM4_3_GP_CalGP21_line3);
nand2 M4_UM4_3_GP_CalGP21_Xo4(M4_UM4_3_GP_CalGP21_line2, M4_UM4_3_GP_CalGP21_line3, M4_UM4_3_Pbus_9);
inv M4_UM4_3_GP_CalGP22_Xo0(M4_Not_XMbus_10, M4_UM4_3_GP_CalGP22_NotA);
inv M4_UM4_3_GP_CalGP22_Xo1(M4_YMbus_10, M4_UM4_3_GP_CalGP22_NotB);
nand2 M4_UM4_3_GP_CalGP22_Xo2(M4_UM4_3_GP_CalGP22_NotA, M4_YMbus_10, M4_UM4_3_GP_CalGP22_line2);
nand2 M4_UM4_3_GP_CalGP22_Xo3(M4_UM4_3_GP_CalGP22_NotB, M4_Not_XMbus_10, M4_UM4_3_GP_CalGP22_line3);
nand2 M4_UM4_3_GP_CalGP22_Xo4(M4_UM4_3_GP_CalGP22_line2, M4_UM4_3_GP_CalGP22_line3, M4_UM4_3_Pbus_10);
inv M4_UM4_3_GP_CalGP23_Xo0(M4_Not_XMbus_11, M4_UM4_3_GP_CalGP23_NotA);
inv M4_UM4_3_GP_CalGP23_Xo1(M4_YMbus_11, M4_UM4_3_GP_CalGP23_NotB);
nand2 M4_UM4_3_GP_CalGP23_Xo2(M4_UM4_3_GP_CalGP23_NotA, M4_YMbus_11, M4_UM4_3_GP_CalGP23_line2);
nand2 M4_UM4_3_GP_CalGP23_Xo3(M4_UM4_3_GP_CalGP23_NotB, M4_Not_XMbus_11, M4_UM4_3_GP_CalGP23_line3);
nand2 M4_UM4_3_GP_CalGP23_Xo4(M4_UM4_3_GP_CalGP23_line2, M4_UM4_3_GP_CalGP23_line3, M4_UM4_3_Pbus_11);
and2 M4_UM4_3_CalcCy_Cla12_0_Cla3_0(M4_UM4_3_Pbus_2, M4_UM4_3_Gbus_1, M4_UM4_3_CalcCy_Cla12_0_line0);
and3 M4_UM4_3_CalcCy_Cla12_0_Cla3_1(M4_UM4_3_Pbus_2, M4_UM4_3_Pbus_1, M4_UM4_3_Gbus_0, M4_UM4_3_CalcCy_Cla12_0_line1);
or3 M4_UM4_3_CalcCy_Cla12_0_Cla3_2(M4_UM4_3_Gbus_2, M4_UM4_3_CalcCy_Cla12_0_line0, M4_UM4_3_CalcCy_Cla12_0_line1, M4_UM4_3_CalcCy_OutCarry2_0);
and2 M4_UM4_3_CalcCy_Cla12_1_Cla5_0(M4_UM4_3_Pbus_7, M4_UM4_3_Gbus_6, M4_UM4_3_CalcCy_Cla12_1_line0);
and3 M4_UM4_3_CalcCy_Cla12_1_Cla5_1(M4_UM4_3_Pbus_7, M4_UM4_3_Pbus_6, M4_UM4_3_Gbus_5, M4_UM4_3_CalcCy_Cla12_1_line1);
and4 M4_UM4_3_CalcCy_Cla12_1_Cla5_2(M4_UM4_3_Pbus_7, M4_UM4_3_Pbus_6, M4_UM4_3_Pbus_5, M4_UM4_3_Gbus_4, M4_UM4_3_CalcCy_Cla12_1_line2);
and5 M4_UM4_3_CalcCy_Cla12_1_Cla5_3(M4_UM4_3_Pbus_7, M4_UM4_3_Pbus_6, M4_UM4_3_Pbus_5, M4_UM4_3_Pbus_4, M4_UM4_3_Gbus_3, M4_UM4_3_CalcCy_Cla12_1_line3);
or5 M4_UM4_3_CalcCy_Cla12_1_Cla5_4(M4_UM4_3_Gbus_7, M4_UM4_3_CalcCy_Cla12_1_line0, M4_UM4_3_CalcCy_Cla12_1_line1, M4_UM4_3_CalcCy_Cla12_1_line2, M4_UM4_3_CalcCy_Cla12_1_line3, M4_UM4_3_CalcCy_OutCarry7_3);
and2 M4_UM4_3_CalcCy_Cla12_2_Cla4_0(M4_UM4_3_Pbus_11, M4_UM4_3_Gbus_10, M4_UM4_3_CalcCy_Cla12_2_line0);
and3 M4_UM4_3_CalcCy_Cla12_2_Cla4_1(M4_UM4_3_Pbus_11, M4_UM4_3_Pbus_10, M4_UM4_3_Gbus_9, M4_UM4_3_CalcCy_Cla12_2_line1);
and4 M4_UM4_3_CalcCy_Cla12_2_Cla4_2(M4_UM4_3_Pbus_11, M4_UM4_3_Pbus_10, M4_UM4_3_Pbus_9, M4_UM4_3_Gbus_8, M4_UM4_3_CalcCy_Cla12_2_line2);
or4 M4_UM4_3_CalcCy_Cla12_2_Cla4_3(M4_UM4_3_Gbus_11, M4_UM4_3_CalcCy_Cla12_2_line0, M4_UM4_3_CalcCy_Cla12_2_line1, M4_UM4_3_CalcCy_Cla12_2_line2, M4_UM4_3_CalcCy_OutCarry11_8);
and5 M4_UM4_3_CalcCy_Cla12_3(M4_UM4_3_Pbus_3, M4_UM4_3_Pbus_4, M4_UM4_3_Pbus_5, M4_UM4_3_Pbus_6, M4_UM4_3_Pbus_7, M4_UM4_3_CalcCy_Prop7_3);
and4 M4_UM4_3_CalcCy_Cla12_4(M4_UM4_3_Pbus_8, M4_UM4_3_Pbus_9, M4_UM4_3_Pbus_10, M4_UM4_3_Pbus_11, M4_UM4_3_CalcCy_Prop11_8);
and2 M4_UM4_3_CalcCy_Cla12_5(M4_UM4_3_CalcCy_Prop7_3, M4_UM4_3_CalcCy_OutCarry2_0, M4_UM4_3_CalcCy_line5);
or2 M4_UM4_3_CalcCy_Cla12_6(M4_UM4_3_CalcCy_OutCarry7_3, M4_UM4_3_CalcCy_line5, M4_UM4_3_CalcCy_OutCarry7_0);
inv M4_UM4_3_CalcCy_Cla12_7(M4_UM4_3_CalcCy_OutCarry7_0, M4_UM4_3_CalcCy_NotOutCarry7_0);
or2 M4_UM4_3_CalcCy_Cla12_8(M4_UM4_3_CalcCy_OutCarry11_8, M4_UM4_3_CalcCy_Prop11_8, M4_UM4_3_CalcCy_line8);
and2 M4_UM4_3_CalcCy_Cla12_9(M4_UM4_3_CalcCy_NotOutCarry7_0, M4_UM4_3_CalcCy_OutCarry11_8, M4_UM4_3_CalcCy_line9);
and2 M4_UM4_3_CalcCy_Cla12_10(M4_UM4_3_CalcCy_line8, M4_UM4_3_CalcCy_OutCarry7_0, M4_UM4_3_CalcCy_line10);
or2 M4_UM4_3_CalcCy_Cla12_11(M4_UM4_3_CalcCy_line9, M4_UM4_3_CalcCy_line10, out329);
and2 M4_UM4_4_GP_CalGP0(M4_Not_XMbus_0, Ybus_0, M4_UM4_4_Gbus_0);
and2 M4_UM4_4_GP_CalGP1(M4_Not_XMbus_1, Ybus_1, M4_UM4_4_Gbus_1);
and2 M4_UM4_4_GP_CalGP2(M4_Not_XMbus_2, Ybus_2, M4_UM4_4_Gbus_2);
and2 M4_UM4_4_GP_CalGP3(M4_Not_XMbus_3, Ybus_3, M4_UM4_4_Gbus_3);
and2 M4_UM4_4_GP_CalGP4(M4_Not_XMbus_4, M4_YMbus_4, M4_UM4_4_Gbus_4);
and2 M4_UM4_4_GP_CalGP5(M4_Not_XMbus_5, M4_YMbus_5, M4_UM4_4_Gbus_5);
and2 M4_UM4_4_GP_CalGP6(M4_Not_XMbus_6, M4_YMbus_6, M4_UM4_4_Gbus_6);
and2 M4_UM4_4_GP_CalGP7(M4_Not_XMbus_7, M4_YMbus_7, M4_UM4_4_Gbus_7);
and2 M4_UM4_4_GP_CalGP8(M4_Not_XMbus_8, M4_YMbus_8, M4_UM4_4_Gbus_8);
and2 M4_UM4_4_GP_CalGP9(M4_Not_XMbus_9, M4_YMbus_9, M4_UM4_4_Gbus_9);
and2 M4_UM4_4_GP_CalGP10(M4_Not_XMbus_10, M4_YMbus_10, M4_UM4_4_Gbus_10);
and2 M4_UM4_4_GP_CalGP11(M4_Not_XMbus_11, M4_YMbus_11, M4_UM4_4_Gbus_11);
inv M4_UM4_4_GP_CalGP12_Xo0(M4_Not_XMbus_0, M4_UM4_4_GP_CalGP12_NotA);
inv M4_UM4_4_GP_CalGP12_Xo1(Ybus_0, M4_UM4_4_GP_CalGP12_NotB);
nand2 M4_UM4_4_GP_CalGP12_Xo2(M4_UM4_4_GP_CalGP12_NotA, Ybus_0, M4_UM4_4_GP_CalGP12_line2);
nand2 M4_UM4_4_GP_CalGP12_Xo3(M4_UM4_4_GP_CalGP12_NotB, M4_Not_XMbus_0, M4_UM4_4_GP_CalGP12_line3);
nand2 M4_UM4_4_GP_CalGP12_Xo4(M4_UM4_4_GP_CalGP12_line2, M4_UM4_4_GP_CalGP12_line3, M4_UM4_4_Pbus_0);
inv M4_UM4_4_GP_CalGP13_Xo0(M4_Not_XMbus_1, M4_UM4_4_GP_CalGP13_NotA);
inv M4_UM4_4_GP_CalGP13_Xo1(Ybus_1, M4_UM4_4_GP_CalGP13_NotB);
nand2 M4_UM4_4_GP_CalGP13_Xo2(M4_UM4_4_GP_CalGP13_NotA, Ybus_1, M4_UM4_4_GP_CalGP13_line2);
nand2 M4_UM4_4_GP_CalGP13_Xo3(M4_UM4_4_GP_CalGP13_NotB, M4_Not_XMbus_1, M4_UM4_4_GP_CalGP13_line3);
nand2 M4_UM4_4_GP_CalGP13_Xo4(M4_UM4_4_GP_CalGP13_line2, M4_UM4_4_GP_CalGP13_line3, M4_UM4_4_Pbus_1);
inv M4_UM4_4_GP_CalGP14_Xo0(M4_Not_XMbus_2, M4_UM4_4_GP_CalGP14_NotA);
inv M4_UM4_4_GP_CalGP14_Xo1(Ybus_2, M4_UM4_4_GP_CalGP14_NotB);
nand2 M4_UM4_4_GP_CalGP14_Xo2(M4_UM4_4_GP_CalGP14_NotA, Ybus_2, M4_UM4_4_GP_CalGP14_line2);
nand2 M4_UM4_4_GP_CalGP14_Xo3(M4_UM4_4_GP_CalGP14_NotB, M4_Not_XMbus_2, M4_UM4_4_GP_CalGP14_line3);
nand2 M4_UM4_4_GP_CalGP14_Xo4(M4_UM4_4_GP_CalGP14_line2, M4_UM4_4_GP_CalGP14_line3, M4_UM4_4_Pbus_2);
inv M4_UM4_4_GP_CalGP15_Xo0(M4_Not_XMbus_3, M4_UM4_4_GP_CalGP15_NotA);
inv M4_UM4_4_GP_CalGP15_Xo1(Ybus_3, M4_UM4_4_GP_CalGP15_NotB);
nand2 M4_UM4_4_GP_CalGP15_Xo2(M4_UM4_4_GP_CalGP15_NotA, Ybus_3, M4_UM4_4_GP_CalGP15_line2);
nand2 M4_UM4_4_GP_CalGP15_Xo3(M4_UM4_4_GP_CalGP15_NotB, M4_Not_XMbus_3, M4_UM4_4_GP_CalGP15_line3);
nand2 M4_UM4_4_GP_CalGP15_Xo4(M4_UM4_4_GP_CalGP15_line2, M4_UM4_4_GP_CalGP15_line3, M4_UM4_4_Pbus_3);
inv M4_UM4_4_GP_CalGP16_Xo0(M4_Not_XMbus_4, M4_UM4_4_GP_CalGP16_NotA);
inv M4_UM4_4_GP_CalGP16_Xo1(M4_YMbus_4, M4_UM4_4_GP_CalGP16_NotB);
nand2 M4_UM4_4_GP_CalGP16_Xo2(M4_UM4_4_GP_CalGP16_NotA, M4_YMbus_4, M4_UM4_4_GP_CalGP16_line2);
nand2 M4_UM4_4_GP_CalGP16_Xo3(M4_UM4_4_GP_CalGP16_NotB, M4_Not_XMbus_4, M4_UM4_4_GP_CalGP16_line3);
nand2 M4_UM4_4_GP_CalGP16_Xo4(M4_UM4_4_GP_CalGP16_line2, M4_UM4_4_GP_CalGP16_line3, M4_UM4_4_Pbus_4);
inv M4_UM4_4_GP_CalGP17_Xo0(M4_Not_XMbus_5, M4_UM4_4_GP_CalGP17_NotA);
inv M4_UM4_4_GP_CalGP17_Xo1(M4_YMbus_5, M4_UM4_4_GP_CalGP17_NotB);
nand2 M4_UM4_4_GP_CalGP17_Xo2(M4_UM4_4_GP_CalGP17_NotA, M4_YMbus_5, M4_UM4_4_GP_CalGP17_line2);
nand2 M4_UM4_4_GP_CalGP17_Xo3(M4_UM4_4_GP_CalGP17_NotB, M4_Not_XMbus_5, M4_UM4_4_GP_CalGP17_line3);
nand2 M4_UM4_4_GP_CalGP17_Xo4(M4_UM4_4_GP_CalGP17_line2, M4_UM4_4_GP_CalGP17_line3, M4_UM4_4_Pbus_5);
inv M4_UM4_4_GP_CalGP18_Xo0(M4_Not_XMbus_6, M4_UM4_4_GP_CalGP18_NotA);
inv M4_UM4_4_GP_CalGP18_Xo1(M4_YMbus_6, M4_UM4_4_GP_CalGP18_NotB);
nand2 M4_UM4_4_GP_CalGP18_Xo2(M4_UM4_4_GP_CalGP18_NotA, M4_YMbus_6, M4_UM4_4_GP_CalGP18_line2);
nand2 M4_UM4_4_GP_CalGP18_Xo3(M4_UM4_4_GP_CalGP18_NotB, M4_Not_XMbus_6, M4_UM4_4_GP_CalGP18_line3);
nand2 M4_UM4_4_GP_CalGP18_Xo4(M4_UM4_4_GP_CalGP18_line2, M4_UM4_4_GP_CalGP18_line3, M4_UM4_4_Pbus_6);
inv M4_UM4_4_GP_CalGP19_Xo0(M4_Not_XMbus_7, M4_UM4_4_GP_CalGP19_NotA);
inv M4_UM4_4_GP_CalGP19_Xo1(M4_YMbus_7, M4_UM4_4_GP_CalGP19_NotB);
nand2 M4_UM4_4_GP_CalGP19_Xo2(M4_UM4_4_GP_CalGP19_NotA, M4_YMbus_7, M4_UM4_4_GP_CalGP19_line2);
nand2 M4_UM4_4_GP_CalGP19_Xo3(M4_UM4_4_GP_CalGP19_NotB, M4_Not_XMbus_7, M4_UM4_4_GP_CalGP19_line3);
nand2 M4_UM4_4_GP_CalGP19_Xo4(M4_UM4_4_GP_CalGP19_line2, M4_UM4_4_GP_CalGP19_line3, M4_UM4_4_Pbus_7);
inv M4_UM4_4_GP_CalGP20_Xo0(M4_Not_XMbus_8, M4_UM4_4_GP_CalGP20_NotA);
inv M4_UM4_4_GP_CalGP20_Xo1(M4_YMbus_8, M4_UM4_4_GP_CalGP20_NotB);
nand2 M4_UM4_4_GP_CalGP20_Xo2(M4_UM4_4_GP_CalGP20_NotA, M4_YMbus_8, M4_UM4_4_GP_CalGP20_line2);
nand2 M4_UM4_4_GP_CalGP20_Xo3(M4_UM4_4_GP_CalGP20_NotB, M4_Not_XMbus_8, M4_UM4_4_GP_CalGP20_line3);
nand2 M4_UM4_4_GP_CalGP20_Xo4(M4_UM4_4_GP_CalGP20_line2, M4_UM4_4_GP_CalGP20_line3, M4_UM4_4_Pbus_8);
inv M4_UM4_4_GP_CalGP21_Xo0(M4_Not_XMbus_9, M4_UM4_4_GP_CalGP21_NotA);
inv M4_UM4_4_GP_CalGP21_Xo1(M4_YMbus_9, M4_UM4_4_GP_CalGP21_NotB);
nand2 M4_UM4_4_GP_CalGP21_Xo2(M4_UM4_4_GP_CalGP21_NotA, M4_YMbus_9, M4_UM4_4_GP_CalGP21_line2);
nand2 M4_UM4_4_GP_CalGP21_Xo3(M4_UM4_4_GP_CalGP21_NotB, M4_Not_XMbus_9, M4_UM4_4_GP_CalGP21_line3);
nand2 M4_UM4_4_GP_CalGP21_Xo4(M4_UM4_4_GP_CalGP21_line2, M4_UM4_4_GP_CalGP21_line3, M4_UM4_4_Pbus_9);
inv M4_UM4_4_GP_CalGP22_Xo0(M4_Not_XMbus_10, M4_UM4_4_GP_CalGP22_NotA);
inv M4_UM4_4_GP_CalGP22_Xo1(M4_YMbus_10, M4_UM4_4_GP_CalGP22_NotB);
nand2 M4_UM4_4_GP_CalGP22_Xo2(M4_UM4_4_GP_CalGP22_NotA, M4_YMbus_10, M4_UM4_4_GP_CalGP22_line2);
nand2 M4_UM4_4_GP_CalGP22_Xo3(M4_UM4_4_GP_CalGP22_NotB, M4_Not_XMbus_10, M4_UM4_4_GP_CalGP22_line3);
nand2 M4_UM4_4_GP_CalGP22_Xo4(M4_UM4_4_GP_CalGP22_line2, M4_UM4_4_GP_CalGP22_line3, M4_UM4_4_Pbus_10);
inv M4_UM4_4_GP_CalGP23_Xo0(M4_Not_XMbus_11, M4_UM4_4_GP_CalGP23_NotA);
inv M4_UM4_4_GP_CalGP23_Xo1(M4_YMbus_11, M4_UM4_4_GP_CalGP23_NotB);
nand2 M4_UM4_4_GP_CalGP23_Xo2(M4_UM4_4_GP_CalGP23_NotA, M4_YMbus_11, M4_UM4_4_GP_CalGP23_line2);
nand2 M4_UM4_4_GP_CalGP23_Xo3(M4_UM4_4_GP_CalGP23_NotB, M4_Not_XMbus_11, M4_UM4_4_GP_CalGP23_line3);
nand2 M4_UM4_4_GP_CalGP23_Xo4(M4_UM4_4_GP_CalGP23_line2, M4_UM4_4_GP_CalGP23_line3, M4_UM4_4_Pbus_11);
and2 M4_UM4_4_CalcCy_Cla12_0_Cla3_0(M4_UM4_4_Pbus_2, M4_UM4_4_Gbus_1, M4_UM4_4_CalcCy_Cla12_0_line0);
and3 M4_UM4_4_CalcCy_Cla12_0_Cla3_1(M4_UM4_4_Pbus_2, M4_UM4_4_Pbus_1, M4_UM4_4_Gbus_0, M4_UM4_4_CalcCy_Cla12_0_line1);
or3 M4_UM4_4_CalcCy_Cla12_0_Cla3_2(M4_UM4_4_Gbus_2, M4_UM4_4_CalcCy_Cla12_0_line0, M4_UM4_4_CalcCy_Cla12_0_line1, M4_UM4_4_CalcCy_OutCarry2_0);
and2 M4_UM4_4_CalcCy_Cla12_1_Cla5_0(M4_UM4_4_Pbus_7, M4_UM4_4_Gbus_6, M4_UM4_4_CalcCy_Cla12_1_line0);
and3 M4_UM4_4_CalcCy_Cla12_1_Cla5_1(M4_UM4_4_Pbus_7, M4_UM4_4_Pbus_6, M4_UM4_4_Gbus_5, M4_UM4_4_CalcCy_Cla12_1_line1);
and4 M4_UM4_4_CalcCy_Cla12_1_Cla5_2(M4_UM4_4_Pbus_7, M4_UM4_4_Pbus_6, M4_UM4_4_Pbus_5, M4_UM4_4_Gbus_4, M4_UM4_4_CalcCy_Cla12_1_line2);
and5 M4_UM4_4_CalcCy_Cla12_1_Cla5_3(M4_UM4_4_Pbus_7, M4_UM4_4_Pbus_6, M4_UM4_4_Pbus_5, M4_UM4_4_Pbus_4, M4_UM4_4_Gbus_3, M4_UM4_4_CalcCy_Cla12_1_line3);
or5 M4_UM4_4_CalcCy_Cla12_1_Cla5_4(M4_UM4_4_Gbus_7, M4_UM4_4_CalcCy_Cla12_1_line0, M4_UM4_4_CalcCy_Cla12_1_line1, M4_UM4_4_CalcCy_Cla12_1_line2, M4_UM4_4_CalcCy_Cla12_1_line3, M4_UM4_4_CalcCy_OutCarry7_3);
and2 M4_UM4_4_CalcCy_Cla12_2_Cla4_0(M4_UM4_4_Pbus_11, M4_UM4_4_Gbus_10, M4_UM4_4_CalcCy_Cla12_2_line0);
and3 M4_UM4_4_CalcCy_Cla12_2_Cla4_1(M4_UM4_4_Pbus_11, M4_UM4_4_Pbus_10, M4_UM4_4_Gbus_9, M4_UM4_4_CalcCy_Cla12_2_line1);
and4 M4_UM4_4_CalcCy_Cla12_2_Cla4_2(M4_UM4_4_Pbus_11, M4_UM4_4_Pbus_10, M4_UM4_4_Pbus_9, M4_UM4_4_Gbus_8, M4_UM4_4_CalcCy_Cla12_2_line2);
or4 M4_UM4_4_CalcCy_Cla12_2_Cla4_3(M4_UM4_4_Gbus_11, M4_UM4_4_CalcCy_Cla12_2_line0, M4_UM4_4_CalcCy_Cla12_2_line1, M4_UM4_4_CalcCy_Cla12_2_line2, M4_UM4_4_CalcCy_OutCarry11_8);
and5 M4_UM4_4_CalcCy_Cla12_3(M4_UM4_4_Pbus_3, M4_UM4_4_Pbus_4, M4_UM4_4_Pbus_5, M4_UM4_4_Pbus_6, M4_UM4_4_Pbus_7, M4_UM4_4_CalcCy_Prop7_3);
and4 M4_UM4_4_CalcCy_Cla12_4(M4_UM4_4_Pbus_8, M4_UM4_4_Pbus_9, M4_UM4_4_Pbus_10, M4_UM4_4_Pbus_11, M4_UM4_4_CalcCy_Prop11_8);
and2 M4_UM4_4_CalcCy_Cla12_5(M4_UM4_4_CalcCy_Prop7_3, M4_UM4_4_CalcCy_OutCarry2_0, M4_UM4_4_CalcCy_line5);
or2 M4_UM4_4_CalcCy_Cla12_6(M4_UM4_4_CalcCy_OutCarry7_3, M4_UM4_4_CalcCy_line5, M4_UM4_4_CalcCy_OutCarry7_0);
inv M4_UM4_4_CalcCy_Cla12_7(M4_UM4_4_CalcCy_OutCarry7_0, M4_UM4_4_CalcCy_NotOutCarry7_0);
or2 M4_UM4_4_CalcCy_Cla12_8(M4_UM4_4_CalcCy_OutCarry11_8, M4_UM4_4_CalcCy_Prop11_8, M4_UM4_4_CalcCy_line8);
and2 M4_UM4_4_CalcCy_Cla12_9(M4_UM4_4_CalcCy_NotOutCarry7_0, M4_UM4_4_CalcCy_OutCarry11_8, M4_UM4_4_CalcCy_line9);
and2 M4_UM4_4_CalcCy_Cla12_10(M4_UM4_4_CalcCy_line8, M4_UM4_4_CalcCy_OutCarry7_0, M4_UM4_4_CalcCy_line10);
or2 M4_UM4_4_CalcCy_Cla12_11(M4_UM4_4_CalcCy_line9, M4_UM4_4_CalcCy_line10, M4_YgX2);
nand2 M4_UM4_5_Xo1_0(out329, M4_YgX2, M4_UM4_5_NotAB);
and2 M4_UM4_5_Xo1_1(out329, M4_UM4_5_NotAB, M4_UM4_5_line1);
and2 M4_UM4_5_Xo1_2(M4_UM4_5_NotAB, M4_YgX2, M4_UM4_5_line2);
or2 M4_UM4_5_Xo1_3(M4_UM4_5_line1, M4_UM4_5_line2, M4_Not_CompCLAs);
inv M4_UM4_6_RIV0(M4_Not_CompCLAs, M4_UM4_6_NotA);
and2 M4_UM4_6_RIV1(M4_Not_CompCLAs, M4_UM4_6_NotA, M4_UM4_6_line1);
or2 M4_UM4_6_RIV2(M4_UM4_6_line1, M4_UM4_6_NotA, CompCLAs);
inv M4_UM4_7(CompCLAs, out231);
inv M5_UM5_0_Inv6_0(in1341, M5_Not_Y1bus_0);
inv M5_UM5_0_Inv6_1(in1348, M5_Not_Y1bus_1);
inv M5_UM5_0_Inv6_2(in1956, M5_Not_Y1bus_2);
inv M5_UM5_0_Inv6_3(in1961, M5_Not_Y1bus_3);
inv M5_UM5_0_Inv6_4(in1966, M5_Not_Y1bus_4);
inv M5_UM5_0_Inv6_5(in1971, M5_Not_Y1bus_5);
inv M5_UM5_1_Inv6_0(in1996, Ybus_10);
inv M5_UM5_1_Inv6_1(in2067, Ybus_11);
inv M5_UM5_1_Inv6_2(in2072, M5_Not_Y2bus_2);
inv M5_UM5_1_Inv6_3(in2078, M5_Not_Y2bus_3);
inv M5_UM5_1_Inv6_4(in2084, M5_Not_Y2bus_4);
inv M5_UM5_1_Inv6_5(in2090, M5_Not_Y2bus_5);
inv M5_UM5_2_Mux6_0_Mux0(ContAlpha, M5_UM5_2_Mux6_0_Not_ContIn);
and2 M5_UM5_2_Mux6_0_Mux1(M5_Not_Y1bus_0, M5_UM5_2_Mux6_0_Not_ContIn, M5_UM5_2_Mux6_0_line1);
and2 M5_UM5_2_Mux6_0_Mux2(Ybus_10, ContAlpha, M5_UM5_2_Mux6_0_line2);
or2 M5_UM5_2_Mux6_0_Mux3(M5_UM5_2_Mux6_0_line1, M5_UM5_2_Mux6_0_line2, Ybus_0);
inv M5_UM5_2_Mux6_1_Mux0(ContAlpha, M5_UM5_2_Mux6_1_Not_ContIn);
and2 M5_UM5_2_Mux6_1_Mux1(M5_Not_Y1bus_1, M5_UM5_2_Mux6_1_Not_ContIn, M5_UM5_2_Mux6_1_line1);
and2 M5_UM5_2_Mux6_1_Mux2(Ybus_11, ContAlpha, M5_UM5_2_Mux6_1_line2);
or2 M5_UM5_2_Mux6_1_Mux3(M5_UM5_2_Mux6_1_line1, M5_UM5_2_Mux6_1_line2, Ybus_1);
inv M5_UM5_2_Mux6_2_Mux0(ContAlpha, M5_UM5_2_Mux6_2_Not_ContIn);
and2 M5_UM5_2_Mux6_2_Mux1(M5_Not_Y1bus_2, M5_UM5_2_Mux6_2_Not_ContIn, M5_UM5_2_Mux6_2_line1);
and2 M5_UM5_2_Mux6_2_Mux2(M5_Not_Y2bus_2, ContAlpha, M5_UM5_2_Mux6_2_line2);
or2 M5_UM5_2_Mux6_2_Mux3(M5_UM5_2_Mux6_2_line1, M5_UM5_2_Mux6_2_line2, Ybus_2);
inv M5_UM5_2_Mux6_3_Mux0(ContAlpha, M5_UM5_2_Mux6_3_Not_ContIn);
and2 M5_UM5_2_Mux6_3_Mux1(M5_Not_Y1bus_3, M5_UM5_2_Mux6_3_Not_ContIn, M5_UM5_2_Mux6_3_line1);
and2 M5_UM5_2_Mux6_3_Mux2(M5_Not_Y2bus_3, ContAlpha, M5_UM5_2_Mux6_3_line2);
or2 M5_UM5_2_Mux6_3_Mux3(M5_UM5_2_Mux6_3_line1, M5_UM5_2_Mux6_3_line2, Ybus_3);
inv M5_UM5_2_Mux6_4_Mux0(ContAlpha, M5_UM5_2_Mux6_4_Not_ContIn);
and2 M5_UM5_2_Mux6_4_Mux1(M5_Not_Y1bus_4, M5_UM5_2_Mux6_4_Not_ContIn, M5_UM5_2_Mux6_4_line1);
and2 M5_UM5_2_Mux6_4_Mux2(M5_Not_Y2bus_4, ContAlpha, M5_UM5_2_Mux6_4_line2);
or2 M5_UM5_2_Mux6_4_Mux3(M5_UM5_2_Mux6_4_line1, M5_UM5_2_Mux6_4_line2, Ybus_4);
inv M5_UM5_2_Mux6_5_Mux0(ContAlpha, M5_UM5_2_Mux6_5_Not_ContIn);
and2 M5_UM5_2_Mux6_5_Mux1(M5_Not_Y1bus_5, M5_UM5_2_Mux6_5_Not_ContIn, M5_UM5_2_Mux6_5_line1);
and2 M5_UM5_2_Mux6_5_Mux2(M5_Not_Y2bus_5, ContAlpha, M5_UM5_2_Mux6_5_line2);
or2 M5_UM5_2_Mux6_5_Mux3(M5_UM5_2_Mux6_5_line1, M5_UM5_2_Mux6_5_line2, Ybus_5);
inv M5_UM5_3_Inv4_0(in1976, Ybus_6);
inv M5_UM5_3_Inv4_1(in1981, Ybus_7);
inv M5_UM5_3_Inv4_2(in1986, Ybus_8);
inv M5_UM5_3_Inv4_3(in1991, Ybus_9);
inv M6_UM6_0_Mux9_0_Mux0(in16, M6_UM6_0_Mux9_0_Not_ContIn);
and2 M6_UM6_0_Mux9_0_Mux1(in19, M6_UM6_0_Mux9_0_Not_ContIn, M6_UM6_0_Mux9_0_line1);
and2 M6_UM6_0_Mux9_0_Mux2(Abus_0, in16, M6_UM6_0_Mux9_0_line2);
or2 M6_UM6_0_Mux9_0_Mux3(M6_UM6_0_Mux9_0_line1, M6_UM6_0_Mux9_0_line2, Zbus_0);
inv M6_UM6_0_Mux9_1_Mux0(in16, M6_UM6_0_Mux9_1_Not_ContIn);
and2 M6_UM6_0_Mux9_1_Mux1(in4, M6_UM6_0_Mux9_1_Not_ContIn, M6_UM6_0_Mux9_1_line1);
and2 M6_UM6_0_Mux9_1_Mux2(Abus_1, in16, M6_UM6_0_Mux9_1_line2);
or2 M6_UM6_0_Mux9_1_Mux3(M6_UM6_0_Mux9_1_line1, M6_UM6_0_Mux9_1_line2, Zbus_1);
inv M6_UM6_0_Mux9_2_Mux0(in16, M6_UM6_0_Mux9_2_Not_ContIn);
and2 M6_UM6_0_Mux9_2_Mux1(in20, M6_UM6_0_Mux9_2_Not_ContIn, M6_UM6_0_Mux9_2_line1);
and2 M6_UM6_0_Mux9_2_Mux2(Abus_2, in16, M6_UM6_0_Mux9_2_line2);
or2 M6_UM6_0_Mux9_2_Mux3(M6_UM6_0_Mux9_2_line1, M6_UM6_0_Mux9_2_line2, Zbus_2);
inv M6_UM6_0_Mux9_3_Mux0(in16, M6_UM6_0_Mux9_3_Not_ContIn);
and2 M6_UM6_0_Mux9_3_Mux1(in5, M6_UM6_0_Mux9_3_Not_ContIn, M6_UM6_0_Mux9_3_line1);
and2 M6_UM6_0_Mux9_3_Mux2(Abus_3, in16, M6_UM6_0_Mux9_3_line2);
or2 M6_UM6_0_Mux9_3_Mux3(M6_UM6_0_Mux9_3_line1, M6_UM6_0_Mux9_3_line2, Zbus_3);
inv M6_UM6_0_Mux9_4_Mux0(in16, M6_UM6_0_Mux9_4_Not_ContIn);
and2 M6_UM6_0_Mux9_4_Mux1(in21, M6_UM6_0_Mux9_4_Not_ContIn, M6_UM6_0_Mux9_4_line1);
and2 M6_UM6_0_Mux9_4_Mux2(Abus_4, in16, M6_UM6_0_Mux9_4_line2);
or2 M6_UM6_0_Mux9_4_Mux3(M6_UM6_0_Mux9_4_line1, M6_UM6_0_Mux9_4_line2, Zbus_4);
inv M6_UM6_0_Mux9_5_Mux0(in16, M6_UM6_0_Mux9_5_Not_ContIn);
and2 M6_UM6_0_Mux9_5_Mux1(in22, M6_UM6_0_Mux9_5_Not_ContIn, M6_UM6_0_Mux9_5_line1);
and2 M6_UM6_0_Mux9_5_Mux2(Abus_5, in16, M6_UM6_0_Mux9_5_line2);
or2 M6_UM6_0_Mux9_5_Mux3(M6_UM6_0_Mux9_5_line1, M6_UM6_0_Mux9_5_line2, Zbus_5);
inv M6_UM6_0_Mux9_6_Mux0(in16, M6_UM6_0_Mux9_6_Not_ContIn);
and2 M6_UM6_0_Mux9_6_Mux1(in23, M6_UM6_0_Mux9_6_Not_ContIn, M6_UM6_0_Mux9_6_line1);
and2 M6_UM6_0_Mux9_6_Mux2(Abus_6, in16, M6_UM6_0_Mux9_6_line2);
or2 M6_UM6_0_Mux9_6_Mux3(M6_UM6_0_Mux9_6_line1, M6_UM6_0_Mux9_6_line2, Zbus_6);
inv M6_UM6_0_Mux9_7_Mux0(in16, M6_UM6_0_Mux9_7_Not_ContIn);
and2 M6_UM6_0_Mux9_7_Mux1(in6, M6_UM6_0_Mux9_7_Not_ContIn, M6_UM6_0_Mux9_7_line1);
and2 M6_UM6_0_Mux9_7_Mux2(Abus_7, in16, M6_UM6_0_Mux9_7_line2);
or2 M6_UM6_0_Mux9_7_Mux3(M6_UM6_0_Mux9_7_line1, M6_UM6_0_Mux9_7_line2, Zbus_7);
inv M6_UM6_0_Mux9_8_Mux0(in16, M6_UM6_0_Mux9_8_Not_ContIn);
and2 M6_UM6_0_Mux9_8_Mux1(in24, M6_UM6_0_Mux9_8_Not_ContIn, M6_UM6_0_Mux9_8_line1);
and2 M6_UM6_0_Mux9_8_Mux2(Abus_8, in16, M6_UM6_0_Mux9_8_line2);
or2 M6_UM6_0_Mux9_8_Mux3(M6_UM6_0_Mux9_8_line1, M6_UM6_0_Mux9_8_line2, Zbus_8);
inv M6_UM6_1_Mux8_0_Mux0(in29, M6_UM6_1_Mux8_0_Not_ContIn);
and2 M6_UM6_1_Mux8_0_Mux1(in25, M6_UM6_1_Mux8_0_Not_ContIn, M6_UM6_1_Mux8_0_line1);
and2 M6_UM6_1_Mux8_0_Mux2(Bbus_0, in29, M6_UM6_1_Mux8_0_line2);
or2 M6_UM6_1_Mux8_0_Mux3(M6_UM6_1_Mux8_0_line1, M6_UM6_1_Mux8_0_line2, Zbus_9);
inv M6_UM6_1_Mux8_1_Mux0(in29, M6_UM6_1_Mux8_1_Not_ContIn);
and2 M6_UM6_1_Mux8_1_Mux1(in32, M6_UM6_1_Mux8_1_Not_ContIn, M6_UM6_1_Mux8_1_line1);
and2 M6_UM6_1_Mux8_1_Mux2(Bbus_1, in29, M6_UM6_1_Mux8_1_line2);
or2 M6_UM6_1_Mux8_1_Mux3(M6_UM6_1_Mux8_1_line1, M6_UM6_1_Mux8_1_line2, Zbus_10);
inv M6_UM6_1_Mux8_2_Mux0(in29, M6_UM6_1_Mux8_2_Not_ContIn);
and2 M6_UM6_1_Mux8_2_Mux1(in26, M6_UM6_1_Mux8_2_Not_ContIn, M6_UM6_1_Mux8_2_line1);
and2 M6_UM6_1_Mux8_2_Mux2(Bbus_2, in29, M6_UM6_1_Mux8_2_line2);
or2 M6_UM6_1_Mux8_2_Mux3(M6_UM6_1_Mux8_2_line1, M6_UM6_1_Mux8_2_line2, Zbus_11);
inv M6_UM6_1_Mux8_3_Mux0(in29, M6_UM6_1_Mux8_3_Not_ContIn);
and2 M6_UM6_1_Mux8_3_Mux1(in33, M6_UM6_1_Mux8_3_Not_ContIn, M6_UM6_1_Mux8_3_line1);
and2 M6_UM6_1_Mux8_3_Mux2(Bbus_3, in29, M6_UM6_1_Mux8_3_line2);
or2 M6_UM6_1_Mux8_3_Mux3(M6_UM6_1_Mux8_3_line1, M6_UM6_1_Mux8_3_line2, Zbus_12);
inv M6_UM6_1_Mux8_4_Mux0(in29, M6_UM6_1_Mux8_4_Not_ContIn);
and2 M6_UM6_1_Mux8_4_Mux1(in27, M6_UM6_1_Mux8_4_Not_ContIn, M6_UM6_1_Mux8_4_line1);
and2 M6_UM6_1_Mux8_4_Mux2(Bbus_4, in29, M6_UM6_1_Mux8_4_line2);
or2 M6_UM6_1_Mux8_4_Mux3(M6_UM6_1_Mux8_4_line1, M6_UM6_1_Mux8_4_line2, Zbus_13);
inv M6_UM6_1_Mux8_5_Mux0(in29, M6_UM6_1_Mux8_5_Not_ContIn);
and2 M6_UM6_1_Mux8_5_Mux1(in34, M6_UM6_1_Mux8_5_Not_ContIn, M6_UM6_1_Mux8_5_line1);
and2 M6_UM6_1_Mux8_5_Mux2(Bbus_5, in29, M6_UM6_1_Mux8_5_line2);
or2 M6_UM6_1_Mux8_5_Mux3(M6_UM6_1_Mux8_5_line1, M6_UM6_1_Mux8_5_line2, Zbus_14);
inv M6_UM6_1_Mux8_6_Mux0(in29, M6_UM6_1_Mux8_6_Not_ContIn);
and2 M6_UM6_1_Mux8_6_Mux1(in35, M6_UM6_1_Mux8_6_Not_ContIn, M6_UM6_1_Mux8_6_line1);
and2 M6_UM6_1_Mux8_6_Mux2(Bbus_6, in29, M6_UM6_1_Mux8_6_line2);
or2 M6_UM6_1_Mux8_6_Mux3(M6_UM6_1_Mux8_6_line1, M6_UM6_1_Mux8_6_line2, Zbus_15);
inv M6_UM6_1_Mux8_7_Mux0(in29, M6_UM6_1_Mux8_7_Not_ContIn);
and2 M6_UM6_1_Mux8_7_Mux1(in28, M6_UM6_1_Mux8_7_Not_ContIn, M6_UM6_1_Mux8_7_line1);
and2 M6_UM6_1_Mux8_7_Mux2(Bbus_7, in29, M6_UM6_1_Mux8_7_line2);
or2 M6_UM6_1_Mux8_7_Mux3(M6_UM6_1_Mux8_7_line1, M6_UM6_1_Mux8_7_line2, Zbus_16);
inv M7_UM7_0_Xr0_Xo0(Zbus_0, M7_UM7_0_Xr0_NotA);
inv M7_UM7_0_Xr0_Xo1(in1341, M7_UM7_0_Xr0_NotB);
nand2 M7_UM7_0_Xr0_Xo2(M7_UM7_0_Xr0_NotA, in1341, M7_UM7_0_Xr0_line2);
nand2 M7_UM7_0_Xr0_Xo3(M7_UM7_0_Xr0_NotB, Zbus_0, M7_UM7_0_Xr0_line3);
nand2 M7_UM7_0_Xr0_Xo4(M7_UM7_0_Xr0_line2, M7_UM7_0_Xr0_line3, M7_XorZW_0);
inv M7_UM7_0_Xr1_Xo0(Zbus_1, M7_UM7_0_Xr1_NotA);
inv M7_UM7_0_Xr1_Xo1(in1348, M7_UM7_0_Xr1_NotB);
nand2 M7_UM7_0_Xr1_Xo2(M7_UM7_0_Xr1_NotA, in1348, M7_UM7_0_Xr1_line2);
nand2 M7_UM7_0_Xr1_Xo3(M7_UM7_0_Xr1_NotB, Zbus_1, M7_UM7_0_Xr1_line3);
nand2 M7_UM7_0_Xr1_Xo4(M7_UM7_0_Xr1_line2, M7_UM7_0_Xr1_line3, M7_XorZW_1);
inv M7_UM7_0_Xr2_Xo0(Zbus_2, M7_UM7_0_Xr2_NotA);
inv M7_UM7_0_Xr2_Xo1(in1956, M7_UM7_0_Xr2_NotB);
nand2 M7_UM7_0_Xr2_Xo2(M7_UM7_0_Xr2_NotA, in1956, M7_UM7_0_Xr2_line2);
nand2 M7_UM7_0_Xr2_Xo3(M7_UM7_0_Xr2_NotB, Zbus_2, M7_UM7_0_Xr2_line3);
nand2 M7_UM7_0_Xr2_Xo4(M7_UM7_0_Xr2_line2, M7_UM7_0_Xr2_line3, M7_XorZW_2);
inv M7_UM7_0_Xr3_Xo0(Zbus_3, M7_UM7_0_Xr3_NotA);
inv M7_UM7_0_Xr3_Xo1(in1961, M7_UM7_0_Xr3_NotB);
nand2 M7_UM7_0_Xr3_Xo2(M7_UM7_0_Xr3_NotA, in1961, M7_UM7_0_Xr3_line2);
nand2 M7_UM7_0_Xr3_Xo3(M7_UM7_0_Xr3_NotB, Zbus_3, M7_UM7_0_Xr3_line3);
nand2 M7_UM7_0_Xr3_Xo4(M7_UM7_0_Xr3_line2, M7_UM7_0_Xr3_line3, M7_XorZW_3);
inv M7_UM7_0_Xr4_Xo0(Zbus_4, M7_UM7_0_Xr4_NotA);
inv M7_UM7_0_Xr4_Xo1(in1966, M7_UM7_0_Xr4_NotB);
nand2 M7_UM7_0_Xr4_Xo2(M7_UM7_0_Xr4_NotA, in1966, M7_UM7_0_Xr4_line2);
nand2 M7_UM7_0_Xr4_Xo3(M7_UM7_0_Xr4_NotB, Zbus_4, M7_UM7_0_Xr4_line3);
nand2 M7_UM7_0_Xr4_Xo4(M7_UM7_0_Xr4_line2, M7_UM7_0_Xr4_line3, M7_XorZW_4);
inv M7_UM7_0_Xr5_Xo0(Zbus_5, M7_UM7_0_Xr5_NotA);
inv M7_UM7_0_Xr5_Xo1(in1971, M7_UM7_0_Xr5_NotB);
nand2 M7_UM7_0_Xr5_Xo2(M7_UM7_0_Xr5_NotA, in1971, M7_UM7_0_Xr5_line2);
nand2 M7_UM7_0_Xr5_Xo3(M7_UM7_0_Xr5_NotB, Zbus_5, M7_UM7_0_Xr5_line3);
nand2 M7_UM7_0_Xr5_Xo4(M7_UM7_0_Xr5_line2, M7_UM7_0_Xr5_line3, M7_XorZW_5);
inv M7_UM7_0_Xr6_Xo0(Zbus_6, M7_UM7_0_Xr6_NotA);
inv M7_UM7_0_Xr6_Xo1(in1976, M7_UM7_0_Xr6_NotB);
nand2 M7_UM7_0_Xr6_Xo2(M7_UM7_0_Xr6_NotA, in1976, M7_UM7_0_Xr6_line2);
nand2 M7_UM7_0_Xr6_Xo3(M7_UM7_0_Xr6_NotB, Zbus_6, M7_UM7_0_Xr6_line3);
nand2 M7_UM7_0_Xr6_Xo4(M7_UM7_0_Xr6_line2, M7_UM7_0_Xr6_line3, M7_XorZW_6);
inv M7_UM7_0_Xr7_Xo0(Zbus_7, M7_UM7_0_Xr7_NotA);
inv M7_UM7_0_Xr7_Xo1(in1981, M7_UM7_0_Xr7_NotB);
nand2 M7_UM7_0_Xr7_Xo2(M7_UM7_0_Xr7_NotA, in1981, M7_UM7_0_Xr7_line2);
nand2 M7_UM7_0_Xr7_Xo3(M7_UM7_0_Xr7_NotB, Zbus_7, M7_UM7_0_Xr7_line3);
nand2 M7_UM7_0_Xr7_Xo4(M7_UM7_0_Xr7_line2, M7_UM7_0_Xr7_line3, M7_XorZW_7);
inv M7_UM7_0_Xr8_Xo0(Zbus_8, M7_UM7_0_Xr8_NotA);
inv M7_UM7_0_Xr8_Xo1(in1986, M7_UM7_0_Xr8_NotB);
nand2 M7_UM7_0_Xr8_Xo2(M7_UM7_0_Xr8_NotA, in1986, M7_UM7_0_Xr8_line2);
nand2 M7_UM7_0_Xr8_Xo3(M7_UM7_0_Xr8_NotB, Zbus_8, M7_UM7_0_Xr8_line3);
nand2 M7_UM7_0_Xr8_Xo4(M7_UM7_0_Xr8_line2, M7_UM7_0_Xr8_line3, M7_XorZW_8);
inv M7_UM7_0_Xr9_Xo0(Zbus_9, M7_UM7_0_Xr9_NotA);
inv M7_UM7_0_Xr9_Xo1(in1991, M7_UM7_0_Xr9_NotB);
nand2 M7_UM7_0_Xr9_Xo2(M7_UM7_0_Xr9_NotA, in1991, M7_UM7_0_Xr9_line2);
nand2 M7_UM7_0_Xr9_Xo3(M7_UM7_0_Xr9_NotB, Zbus_9, M7_UM7_0_Xr9_line3);
nand2 M7_UM7_0_Xr9_Xo4(M7_UM7_0_Xr9_line2, M7_UM7_0_Xr9_line3, M7_XorZW_9);
inv M7_UM7_0_Xr10_Xo0(Zbus_10, M7_UM7_0_Xr10_NotA);
inv M7_UM7_0_Xr10_Xo1(in1996, M7_UM7_0_Xr10_NotB);
nand2 M7_UM7_0_Xr10_Xo2(M7_UM7_0_Xr10_NotA, in1996, M7_UM7_0_Xr10_line2);
nand2 M7_UM7_0_Xr10_Xo3(M7_UM7_0_Xr10_NotB, Zbus_10, M7_UM7_0_Xr10_line3);
nand2 M7_UM7_0_Xr10_Xo4(M7_UM7_0_Xr10_line2, M7_UM7_0_Xr10_line3, M7_XorZW_10);
inv M7_UM7_0_Xr11_Xo0(Zbus_11, M7_UM7_0_Xr11_NotA);
inv M7_UM7_0_Xr11_Xo1(in2067, M7_UM7_0_Xr11_NotB);
nand2 M7_UM7_0_Xr11_Xo2(M7_UM7_0_Xr11_NotA, in2067, M7_UM7_0_Xr11_line2);
nand2 M7_UM7_0_Xr11_Xo3(M7_UM7_0_Xr11_NotB, Zbus_11, M7_UM7_0_Xr11_line3);
nand2 M7_UM7_0_Xr11_Xo4(M7_UM7_0_Xr11_line2, M7_UM7_0_Xr11_line3, M7_XorZW_11);
inv M7_UM7_0_Xr12_Xo0(Zbus_12, M7_UM7_0_Xr12_NotA);
inv M7_UM7_0_Xr12_Xo1(in2072, M7_UM7_0_Xr12_NotB);
nand2 M7_UM7_0_Xr12_Xo2(M7_UM7_0_Xr12_NotA, in2072, M7_UM7_0_Xr12_line2);
nand2 M7_UM7_0_Xr12_Xo3(M7_UM7_0_Xr12_NotB, Zbus_12, M7_UM7_0_Xr12_line3);
nand2 M7_UM7_0_Xr12_Xo4(M7_UM7_0_Xr12_line2, M7_UM7_0_Xr12_line3, M7_XorZW_12);
inv M7_UM7_0_Xr13_Xo0(Zbus_13, M7_UM7_0_Xr13_NotA);
inv M7_UM7_0_Xr13_Xo1(in2078, M7_UM7_0_Xr13_NotB);
nand2 M7_UM7_0_Xr13_Xo2(M7_UM7_0_Xr13_NotA, in2078, M7_UM7_0_Xr13_line2);
nand2 M7_UM7_0_Xr13_Xo3(M7_UM7_0_Xr13_NotB, Zbus_13, M7_UM7_0_Xr13_line3);
nand2 M7_UM7_0_Xr13_Xo4(M7_UM7_0_Xr13_line2, M7_UM7_0_Xr13_line3, M7_XorZW_13);
inv M7_UM7_0_Xr14_Xo0(Zbus_14, M7_UM7_0_Xr14_NotA);
inv M7_UM7_0_Xr14_Xo1(in2084, M7_UM7_0_Xr14_NotB);
nand2 M7_UM7_0_Xr14_Xo2(M7_UM7_0_Xr14_NotA, in2084, M7_UM7_0_Xr14_line2);
nand2 M7_UM7_0_Xr14_Xo3(M7_UM7_0_Xr14_NotB, Zbus_14, M7_UM7_0_Xr14_line3);
nand2 M7_UM7_0_Xr14_Xo4(M7_UM7_0_Xr14_line2, M7_UM7_0_Xr14_line3, M7_XorZW_14);
inv M7_UM7_0_Xr15_Xo0(Zbus_15, M7_UM7_0_Xr15_NotA);
inv M7_UM7_0_Xr15_Xo1(in2090, M7_UM7_0_Xr15_NotB);
nand2 M7_UM7_0_Xr15_Xo2(M7_UM7_0_Xr15_NotA, in2090, M7_UM7_0_Xr15_line2);
nand2 M7_UM7_0_Xr15_Xo3(M7_UM7_0_Xr15_NotB, Zbus_15, M7_UM7_0_Xr15_line3);
nand2 M7_UM7_0_Xr15_Xo4(M7_UM7_0_Xr15_line2, M7_UM7_0_Xr15_line3, M7_XorZW_15);
inv M7_UM7_0_Xr16_Xo0(Zbus_16, M7_UM7_0_Xr16_NotA);
inv M7_UM7_0_Xr16_Xo1(gnd, M7_UM7_0_Xr16_NotB);
nand2 M7_UM7_0_Xr16_Xo2(M7_UM7_0_Xr16_NotA, gnd, M7_UM7_0_Xr16_line2);
nand2 M7_UM7_0_Xr16_Xo3(M7_UM7_0_Xr16_NotB, Zbus_16, M7_UM7_0_Xr16_line3);
nand2 M7_UM7_0_Xr16_Xo4(M7_UM7_0_Xr16_line2, M7_UM7_0_Xr16_line3, M7_XorZW_16);
and5 M7_UM7_1_A0(M7_XorZW_0, M7_XorZW_1, M7_XorZW_2, M7_XorZW_3, M7_XorZW_4, M7_UM7_1_line0);
and5 M7_UM7_1_A1(M7_XorZW_5, M7_XorZW_6, M7_XorZW_7, M7_XorZW_8, M7_XorZW_9, M7_UM7_1_line1);
and2 M7_UM7_1_A2(M7_UM7_1_line0, M7_UM7_1_line1, M7_UM7_1_line2);
and2 M7_UM7_1_A3(M7_XorZW_10, M7_XorZW_11, M7_UM7_1_line3);
and5 M7_UM7_1_A4(M7_XorZW_12, M7_XorZW_13, M7_XorZW_14, M7_XorZW_15, M7_XorZW_16, M7_UM7_1_line4);
and2 M7_UM7_1_A5(M7_UM7_1_line3, M7_UM7_1_line4, M7_UM7_1_line5);
and3 M7_UM7_1_A6(M7_UM7_1_line2, M7_UM7_1_line5, in11, out311);
inv M7_UM7_2(out311, out150);
and4 M8_UM8_0_SCL0(in44, in132, in82, in96, M8_UM8_0_line0);
and4 M8_UM8_0_SCL1(in69, in120, in57, in108, M8_UM8_0_line1);
and2 M8_UM8_0_SCL2(M8_UM8_0_line0, M8_UM8_0_line1, out325);
inv M8_UM8_0_SCL3(out325, out261);
inv M8_UM8_0_SCL4(in2106, M8_UM8_0_NotPar2);
inv M8_UM8_0_SCL5(in567, M8_UM8_0_NotPar3);
or2 M8_UM8_0_SCL6(M8_UM8_0_NotPar2, M8_UM8_0_line0, M8_UM8_0_line6);
or2 M8_UM8_0_SCL7(M8_UM8_0_NotPar3, M8_UM8_0_line1, M8_UM8_0_line7);
and2 M8_UM8_0_SCL8(M8_UM8_0_line6, M8_UM8_0_line7, out319);
inv M8_UM8_0_SCL9(in44, out218);
inv M8_UM8_0_SCL10(in132, out219);
inv M8_UM8_0_SCL11(in82, out220);
inv M8_UM8_0_SCL12(in96, out221);
inv M8_UM8_0_SCL13(in69, out235);
inv M8_UM8_0_SCL14(in120, out236);
inv M8_UM8_0_SCL15(in57, out237);
inv M8_UM8_0_SCL16(in108, out238);
inv M8_UM8_1_PT0_Xo0(Abus_0, M8_UM8_1_PT0_NotA);
inv M8_UM8_1_PT0_Xo1(Abus_1, M8_UM8_1_PT0_NotB);
nand2 M8_UM8_1_PT0_Xo2(M8_UM8_1_PT0_NotA, Abus_1, M8_UM8_1_PT0_line2);
nand2 M8_UM8_1_PT0_Xo3(M8_UM8_1_PT0_NotB, Abus_0, M8_UM8_1_PT0_line3);
nand2 M8_UM8_1_PT0_Xo4(M8_UM8_1_PT0_line2, M8_UM8_1_PT0_line3, M8_UM8_1_line0);
inv M8_UM8_1_PT1_Xo0(Abus_2, M8_UM8_1_PT1_NotA);
inv M8_UM8_1_PT1_Xo1(Abus_3, M8_UM8_1_PT1_NotB);
nand2 M8_UM8_1_PT1_Xo2(M8_UM8_1_PT1_NotA, Abus_3, M8_UM8_1_PT1_line2);
nand2 M8_UM8_1_PT1_Xo3(M8_UM8_1_PT1_NotB, Abus_2, M8_UM8_1_PT1_line3);
nand2 M8_UM8_1_PT1_Xo4(M8_UM8_1_PT1_line2, M8_UM8_1_PT1_line3, M8_UM8_1_line1);
inv M8_UM8_1_PT2_Xo0(Abus_4, M8_UM8_1_PT2_NotA);
inv M8_UM8_1_PT2_Xo1(Abus_5, M8_UM8_1_PT2_NotB);
nand2 M8_UM8_1_PT2_Xo2(M8_UM8_1_PT2_NotA, Abus_5, M8_UM8_1_PT2_line2);
nand2 M8_UM8_1_PT2_Xo3(M8_UM8_1_PT2_NotB, Abus_4, M8_UM8_1_PT2_line3);
nand2 M8_UM8_1_PT2_Xo4(M8_UM8_1_PT2_line2, M8_UM8_1_PT2_line3, M8_UM8_1_line2);
inv M8_UM8_1_PT3_Xo0(Abus_6, M8_UM8_1_PT3_NotA);
inv M8_UM8_1_PT3_Xo1(Abus_7, M8_UM8_1_PT3_NotB);
nand2 M8_UM8_1_PT3_Xo2(M8_UM8_1_PT3_NotA, Abus_7, M8_UM8_1_PT3_line2);
nand2 M8_UM8_1_PT3_Xo3(M8_UM8_1_PT3_NotB, Abus_6, M8_UM8_1_PT3_line3);
nand2 M8_UM8_1_PT3_Xo4(M8_UM8_1_PT3_line2, M8_UM8_1_PT3_line3, M8_UM8_1_line3);
inv M8_UM8_1_PT4_Xo0(Abus_8, M8_UM8_1_PT4_NotA);
inv M8_UM8_1_PT4_Xo1(Abus_9, M8_UM8_1_PT4_NotB);
nand2 M8_UM8_1_PT4_Xo2(M8_UM8_1_PT4_NotA, Abus_9, M8_UM8_1_PT4_line2);
nand2 M8_UM8_1_PT4_Xo3(M8_UM8_1_PT4_NotB, Abus_8, M8_UM8_1_PT4_line3);
nand2 M8_UM8_1_PT4_Xo4(M8_UM8_1_PT4_line2, M8_UM8_1_PT4_line3, M8_UM8_1_line4);
inv M8_UM8_1_PT5_Xo3_0(M8_UM8_1_line0, M8_UM8_1_PT5_NotA);
inv M8_UM8_1_PT5_Xo3_1(M8_UM8_1_line1, M8_UM8_1_PT5_NotB);
inv M8_UM8_1_PT5_Xo3_2(M8_UM8_1_line2, M8_UM8_1_PT5_NotC);
and3 M8_UM8_1_PT5_Xo3_3(M8_UM8_1_PT5_NotA, M8_UM8_1_PT5_NotB, M8_UM8_1_line2, M8_UM8_1_PT5_line3);
and3 M8_UM8_1_PT5_Xo3_4(M8_UM8_1_PT5_NotA, M8_UM8_1_line1, M8_UM8_1_PT5_NotC, M8_UM8_1_PT5_line4);
and3 M8_UM8_1_PT5_Xo3_5(M8_UM8_1_line0, M8_UM8_1_PT5_NotB, M8_UM8_1_PT5_NotC, M8_UM8_1_PT5_line5);
and3 M8_UM8_1_PT5_Xo3_6(M8_UM8_1_line0, M8_UM8_1_line1, M8_UM8_1_line2, M8_UM8_1_PT5_line6);
nor2 M8_UM8_1_PT5_Xo3_7(M8_UM8_1_PT5_line3, M8_UM8_1_PT5_line4, M8_UM8_1_PT5_line7);
nor2 M8_UM8_1_PT5_Xo3_8(M8_UM8_1_PT5_line5, M8_UM8_1_PT5_line6, M8_UM8_1_PT5_line8);
nand2 M8_UM8_1_PT5_Xo3_9(M8_UM8_1_PT5_line7, M8_UM8_1_PT5_line8, M8_UM8_1_line5);
inv M8_UM8_1_PT6_Xo0(M8_UM8_1_line3, M8_UM8_1_PT6_NotA);
inv M8_UM8_1_PT6_Xo1(M8_UM8_1_line4, M8_UM8_1_PT6_NotB);
nand2 M8_UM8_1_PT6_Xo2(M8_UM8_1_PT6_NotA, M8_UM8_1_line4, M8_UM8_1_PT6_line2);
nand2 M8_UM8_1_PT6_Xo3(M8_UM8_1_PT6_NotB, M8_UM8_1_line3, M8_UM8_1_PT6_line3);
nand2 M8_UM8_1_PT6_Xo4(M8_UM8_1_PT6_line2, M8_UM8_1_PT6_line3, M8_UM8_1_line6);
inv M8_UM8_1_PT7_Xo0(M8_UM8_1_line5, M8_UM8_1_PT7_NotA);
inv M8_UM8_1_PT7_Xo1(M8_UM8_1_line6, M8_UM8_1_PT7_NotB);
nand2 M8_UM8_1_PT7_Xo2(M8_UM8_1_PT7_NotA, M8_UM8_1_line6, M8_UM8_1_PT7_line2);
nand2 M8_UM8_1_PT7_Xo3(M8_UM8_1_PT7_NotB, M8_UM8_1_line5, M8_UM8_1_PT7_line3);
nand2 M8_UM8_1_PT7_Xo4(M8_UM8_1_PT7_line2, M8_UM8_1_PT7_line3, M8_ParA);
inv M8_UM8_2_PT0_Xo0(Bbus_0, M8_UM8_2_PT0_NotA);
inv M8_UM8_2_PT0_Xo1(Bbus_1, M8_UM8_2_PT0_NotB);
nand2 M8_UM8_2_PT0_Xo2(M8_UM8_2_PT0_NotA, Bbus_1, M8_UM8_2_PT0_line2);
nand2 M8_UM8_2_PT0_Xo3(M8_UM8_2_PT0_NotB, Bbus_0, M8_UM8_2_PT0_line3);
nand2 M8_UM8_2_PT0_Xo4(M8_UM8_2_PT0_line2, M8_UM8_2_PT0_line3, M8_UM8_2_line0);
inv M8_UM8_2_PT1_Xo0(Bbus_2, M8_UM8_2_PT1_NotA);
inv M8_UM8_2_PT1_Xo1(Bbus_3, M8_UM8_2_PT1_NotB);
nand2 M8_UM8_2_PT1_Xo2(M8_UM8_2_PT1_NotA, Bbus_3, M8_UM8_2_PT1_line2);
nand2 M8_UM8_2_PT1_Xo3(M8_UM8_2_PT1_NotB, Bbus_2, M8_UM8_2_PT1_line3);
nand2 M8_UM8_2_PT1_Xo4(M8_UM8_2_PT1_line2, M8_UM8_2_PT1_line3, M8_UM8_2_line1);
inv M8_UM8_2_PT2_Xo0(Bbus_4, M8_UM8_2_PT2_NotA);
inv M8_UM8_2_PT2_Xo1(Bbus_5, M8_UM8_2_PT2_NotB);
nand2 M8_UM8_2_PT2_Xo2(M8_UM8_2_PT2_NotA, Bbus_5, M8_UM8_2_PT2_line2);
nand2 M8_UM8_2_PT2_Xo3(M8_UM8_2_PT2_NotB, Bbus_4, M8_UM8_2_PT2_line3);
nand2 M8_UM8_2_PT2_Xo4(M8_UM8_2_PT2_line2, M8_UM8_2_PT2_line3, M8_UM8_2_line2);
inv M8_UM8_2_PT3_Xo0(Bbus_6, M8_UM8_2_PT3_NotA);
inv M8_UM8_2_PT3_Xo1(Bbus_7, M8_UM8_2_PT3_NotB);
nand2 M8_UM8_2_PT3_Xo2(M8_UM8_2_PT3_NotA, Bbus_7, M8_UM8_2_PT3_line2);
nand2 M8_UM8_2_PT3_Xo3(M8_UM8_2_PT3_NotB, Bbus_6, M8_UM8_2_PT3_line3);
nand2 M8_UM8_2_PT3_Xo4(M8_UM8_2_PT3_line2, M8_UM8_2_PT3_line3, M8_UM8_2_line3);
inv M8_UM8_2_PT4_Xo0(Bbus_8, M8_UM8_2_PT4_NotA);
inv M8_UM8_2_PT4_Xo1(Bbus_9, M8_UM8_2_PT4_NotB);
nand2 M8_UM8_2_PT4_Xo2(M8_UM8_2_PT4_NotA, Bbus_9, M8_UM8_2_PT4_line2);
nand2 M8_UM8_2_PT4_Xo3(M8_UM8_2_PT4_NotB, Bbus_8, M8_UM8_2_PT4_line3);
nand2 M8_UM8_2_PT4_Xo4(M8_UM8_2_PT4_line2, M8_UM8_2_PT4_line3, M8_UM8_2_line4);
inv M8_UM8_2_PT5_Xo3_0(M8_UM8_2_line0, M8_UM8_2_PT5_NotA);
inv M8_UM8_2_PT5_Xo3_1(M8_UM8_2_line1, M8_UM8_2_PT5_NotB);
inv M8_UM8_2_PT5_Xo3_2(M8_UM8_2_line2, M8_UM8_2_PT5_NotC);
and3 M8_UM8_2_PT5_Xo3_3(M8_UM8_2_PT5_NotA, M8_UM8_2_PT5_NotB, M8_UM8_2_line2, M8_UM8_2_PT5_line3);
and3 M8_UM8_2_PT5_Xo3_4(M8_UM8_2_PT5_NotA, M8_UM8_2_line1, M8_UM8_2_PT5_NotC, M8_UM8_2_PT5_line4);
and3 M8_UM8_2_PT5_Xo3_5(M8_UM8_2_line0, M8_UM8_2_PT5_NotB, M8_UM8_2_PT5_NotC, M8_UM8_2_PT5_line5);
and3 M8_UM8_2_PT5_Xo3_6(M8_UM8_2_line0, M8_UM8_2_line1, M8_UM8_2_line2, M8_UM8_2_PT5_line6);
nor2 M8_UM8_2_PT5_Xo3_7(M8_UM8_2_PT5_line3, M8_UM8_2_PT5_line4, M8_UM8_2_PT5_line7);
nor2 M8_UM8_2_PT5_Xo3_8(M8_UM8_2_PT5_line5, M8_UM8_2_PT5_line6, M8_UM8_2_PT5_line8);
nand2 M8_UM8_2_PT5_Xo3_9(M8_UM8_2_PT5_line7, M8_UM8_2_PT5_line8, M8_UM8_2_line5);
inv M8_UM8_2_PT6_Xo0(M8_UM8_2_line3, M8_UM8_2_PT6_NotA);
inv M8_UM8_2_PT6_Xo1(M8_UM8_2_line4, M8_UM8_2_PT6_NotB);
nand2 M8_UM8_2_PT6_Xo2(M8_UM8_2_PT6_NotA, M8_UM8_2_line4, M8_UM8_2_PT6_line2);
nand2 M8_UM8_2_PT6_Xo3(M8_UM8_2_PT6_NotB, M8_UM8_2_line3, M8_UM8_2_PT6_line3);
nand2 M8_UM8_2_PT6_Xo4(M8_UM8_2_PT6_line2, M8_UM8_2_PT6_line3, M8_UM8_2_line6);
inv M8_UM8_2_PT7_Xo0(M8_UM8_2_line5, M8_UM8_2_PT7_NotA);
inv M8_UM8_2_PT7_Xo1(M8_UM8_2_line6, M8_UM8_2_PT7_NotB);
nand2 M8_UM8_2_PT7_Xo2(M8_UM8_2_PT7_NotA, M8_UM8_2_line6, M8_UM8_2_PT7_line2);
nand2 M8_UM8_2_PT7_Xo3(M8_UM8_2_PT7_NotB, M8_UM8_2_line5, M8_UM8_2_PT7_line3);
nand2 M8_UM8_2_PT7_Xo4(M8_UM8_2_PT7_line2, M8_UM8_2_PT7_line3, M8_ParB);
inv M8_UM8_3_PT0_Xo0(in1956, M8_UM8_3_PT0_NotA);
inv M8_UM8_3_PT0_Xo1(in1961, M8_UM8_3_PT0_NotB);
nand2 M8_UM8_3_PT0_Xo2(M8_UM8_3_PT0_NotA, in1961, M8_UM8_3_PT0_line2);
nand2 M8_UM8_3_PT0_Xo3(M8_UM8_3_PT0_NotB, in1956, M8_UM8_3_PT0_line3);
nand2 M8_UM8_3_PT0_Xo4(M8_UM8_3_PT0_line2, M8_UM8_3_PT0_line3, M8_UM8_3_line0);
inv M8_UM8_3_PT1_Xo0(in1966, M8_UM8_3_PT1_NotA);
inv M8_UM8_3_PT1_Xo1(in1971, M8_UM8_3_PT1_NotB);
nand2 M8_UM8_3_PT1_Xo2(M8_UM8_3_PT1_NotA, in1971, M8_UM8_3_PT1_line2);
nand2 M8_UM8_3_PT1_Xo3(M8_UM8_3_PT1_NotB, in1966, M8_UM8_3_PT1_line3);
nand2 M8_UM8_3_PT1_Xo4(M8_UM8_3_PT1_line2, M8_UM8_3_PT1_line3, M8_UM8_3_line1);
inv M8_UM8_3_PT2_Xo0(in1976, M8_UM8_3_PT2_NotA);
inv M8_UM8_3_PT2_Xo1(in1981, M8_UM8_3_PT2_NotB);
nand2 M8_UM8_3_PT2_Xo2(M8_UM8_3_PT2_NotA, in1981, M8_UM8_3_PT2_line2);
nand2 M8_UM8_3_PT2_Xo3(M8_UM8_3_PT2_NotB, in1976, M8_UM8_3_PT2_line3);
nand2 M8_UM8_3_PT2_Xo4(M8_UM8_3_PT2_line2, M8_UM8_3_PT2_line3, M8_UM8_3_line2);
inv M8_UM8_3_PT3_Xo0(in1986, M8_UM8_3_PT3_NotA);
inv M8_UM8_3_PT3_Xo1(in1991, M8_UM8_3_PT3_NotB);
nand2 M8_UM8_3_PT3_Xo2(M8_UM8_3_PT3_NotA, in1991, M8_UM8_3_PT3_line2);
nand2 M8_UM8_3_PT3_Xo3(M8_UM8_3_PT3_NotB, in1986, M8_UM8_3_PT3_line3);
nand2 M8_UM8_3_PT3_Xo4(M8_UM8_3_PT3_line2, M8_UM8_3_PT3_line3, M8_UM8_3_line3);
inv M8_UM8_3_PT4_Xo0(in1996, M8_UM8_3_PT4_NotA);
inv M8_UM8_3_PT4_Xo1(in2474, M8_UM8_3_PT4_NotB);
nand2 M8_UM8_3_PT4_Xo2(M8_UM8_3_PT4_NotA, in2474, M8_UM8_3_PT4_line2);
nand2 M8_UM8_3_PT4_Xo3(M8_UM8_3_PT4_NotB, in1996, M8_UM8_3_PT4_line3);
nand2 M8_UM8_3_PT4_Xo4(M8_UM8_3_PT4_line2, M8_UM8_3_PT4_line3, M8_UM8_3_line4);
inv M8_UM8_3_PT5_Xo3_0(M8_UM8_3_line0, M8_UM8_3_PT5_NotA);
inv M8_UM8_3_PT5_Xo3_1(M8_UM8_3_line1, M8_UM8_3_PT5_NotB);
inv M8_UM8_3_PT5_Xo3_2(M8_UM8_3_line2, M8_UM8_3_PT5_NotC);
and3 M8_UM8_3_PT5_Xo3_3(M8_UM8_3_PT5_NotA, M8_UM8_3_PT5_NotB, M8_UM8_3_line2, M8_UM8_3_PT5_line3);
and3 M8_UM8_3_PT5_Xo3_4(M8_UM8_3_PT5_NotA, M8_UM8_3_line1, M8_UM8_3_PT5_NotC, M8_UM8_3_PT5_line4);
and3 M8_UM8_3_PT5_Xo3_5(M8_UM8_3_line0, M8_UM8_3_PT5_NotB, M8_UM8_3_PT5_NotC, M8_UM8_3_PT5_line5);
and3 M8_UM8_3_PT5_Xo3_6(M8_UM8_3_line0, M8_UM8_3_line1, M8_UM8_3_line2, M8_UM8_3_PT5_line6);
nor2 M8_UM8_3_PT5_Xo3_7(M8_UM8_3_PT5_line3, M8_UM8_3_PT5_line4, M8_UM8_3_PT5_line7);
nor2 M8_UM8_3_PT5_Xo3_8(M8_UM8_3_PT5_line5, M8_UM8_3_PT5_line6, M8_UM8_3_PT5_line8);
nand2 M8_UM8_3_PT5_Xo3_9(M8_UM8_3_PT5_line7, M8_UM8_3_PT5_line8, M8_UM8_3_line5);
inv M8_UM8_3_PT6_Xo0(M8_UM8_3_line3, M8_UM8_3_PT6_NotA);
inv M8_UM8_3_PT6_Xo1(M8_UM8_3_line4, M8_UM8_3_PT6_NotB);
nand2 M8_UM8_3_PT6_Xo2(M8_UM8_3_PT6_NotA, M8_UM8_3_line4, M8_UM8_3_PT6_line2);
nand2 M8_UM8_3_PT6_Xo3(M8_UM8_3_PT6_NotB, M8_UM8_3_line3, M8_UM8_3_PT6_line3);
nand2 M8_UM8_3_PT6_Xo4(M8_UM8_3_PT6_line2, M8_UM8_3_PT6_line3, M8_UM8_3_line6);
inv M8_UM8_3_PT7_Xo0(M8_UM8_3_line5, M8_UM8_3_PT7_NotA);
inv M8_UM8_3_PT7_Xo1(M8_UM8_3_line6, M8_UM8_3_PT7_NotB);
nand2 M8_UM8_3_PT7_Xo2(M8_UM8_3_PT7_NotA, M8_UM8_3_line6, M8_UM8_3_PT7_line2);
nand2 M8_UM8_3_PT7_Xo3(M8_UM8_3_PT7_NotB, M8_UM8_3_line5, M8_UM8_3_PT7_line3);
nand2 M8_UM8_3_PT7_Xo4(M8_UM8_3_PT7_line2, M8_UM8_3_PT7_line3, M8_ParQ);
inv M8_UM8_4_PT0_Xo0(in1341, M8_UM8_4_PT0_NotA);
inv M8_UM8_4_PT0_Xo1(in1348, M8_UM8_4_PT0_NotB);
nand2 M8_UM8_4_PT0_Xo2(M8_UM8_4_PT0_NotA, in1348, M8_UM8_4_PT0_line2);
nand2 M8_UM8_4_PT0_Xo3(M8_UM8_4_PT0_NotB, in1341, M8_UM8_4_PT0_line3);
nand2 M8_UM8_4_PT0_Xo4(M8_UM8_4_PT0_line2, M8_UM8_4_PT0_line3, M8_UM8_4_line0);
inv M8_UM8_4_PT1_Xo0(in2427, M8_UM8_4_PT1_NotA);
inv M8_UM8_4_PT1_Xo1(in2430, M8_UM8_4_PT1_NotB);
nand2 M8_UM8_4_PT1_Xo2(M8_UM8_4_PT1_NotA, in2430, M8_UM8_4_PT1_line2);
nand2 M8_UM8_4_PT1_Xo3(M8_UM8_4_PT1_NotB, in2427, M8_UM8_4_PT1_line3);
nand2 M8_UM8_4_PT1_Xo4(M8_UM8_4_PT1_line2, M8_UM8_4_PT1_line3, M8_UM8_4_line1);
inv M8_UM8_4_PT2_Xo0(in2435, M8_UM8_4_PT2_NotA);
inv M8_UM8_4_PT2_Xo1(in2438, M8_UM8_4_PT2_NotB);
nand2 M8_UM8_4_PT2_Xo2(M8_UM8_4_PT2_NotA, in2438, M8_UM8_4_PT2_line2);
nand2 M8_UM8_4_PT2_Xo3(M8_UM8_4_PT2_NotB, in2435, M8_UM8_4_PT2_line3);
nand2 M8_UM8_4_PT2_Xo4(M8_UM8_4_PT2_line2, M8_UM8_4_PT2_line3, M8_UM8_4_line2);
inv M8_UM8_4_PT3_Xo0(in2443, M8_UM8_4_PT3_NotA);
inv M8_UM8_4_PT3_Xo1(in2446, M8_UM8_4_PT3_NotB);
nand2 M8_UM8_4_PT3_Xo2(M8_UM8_4_PT3_NotA, in2446, M8_UM8_4_PT3_line2);
nand2 M8_UM8_4_PT3_Xo3(M8_UM8_4_PT3_NotB, in2443, M8_UM8_4_PT3_line3);
nand2 M8_UM8_4_PT3_Xo4(M8_UM8_4_PT3_line2, M8_UM8_4_PT3_line3, M8_UM8_4_line3);
inv M8_UM8_4_PT4_Xo0(in2451, M8_UM8_4_PT4_NotA);
inv M8_UM8_4_PT4_Xo1(in2454, M8_UM8_4_PT4_NotB);
nand2 M8_UM8_4_PT4_Xo2(M8_UM8_4_PT4_NotA, in2454, M8_UM8_4_PT4_line2);
nand2 M8_UM8_4_PT4_Xo3(M8_UM8_4_PT4_NotB, in2451, M8_UM8_4_PT4_line3);
nand2 M8_UM8_4_PT4_Xo4(M8_UM8_4_PT4_line2, M8_UM8_4_PT4_line3, M8_UM8_4_line4);
inv M8_UM8_4_PT5_Xo3_0(M8_UM8_4_line0, M8_UM8_4_PT5_NotA);
inv M8_UM8_4_PT5_Xo3_1(M8_UM8_4_line1, M8_UM8_4_PT5_NotB);
inv M8_UM8_4_PT5_Xo3_2(M8_UM8_4_line2, M8_UM8_4_PT5_NotC);
and3 M8_UM8_4_PT5_Xo3_3(M8_UM8_4_PT5_NotA, M8_UM8_4_PT5_NotB, M8_UM8_4_line2, M8_UM8_4_PT5_line3);
and3 M8_UM8_4_PT5_Xo3_4(M8_UM8_4_PT5_NotA, M8_UM8_4_line1, M8_UM8_4_PT5_NotC, M8_UM8_4_PT5_line4);
and3 M8_UM8_4_PT5_Xo3_5(M8_UM8_4_line0, M8_UM8_4_PT5_NotB, M8_UM8_4_PT5_NotC, M8_UM8_4_PT5_line5);
and3 M8_UM8_4_PT5_Xo3_6(M8_UM8_4_line0, M8_UM8_4_line1, M8_UM8_4_line2, M8_UM8_4_PT5_line6);
nor2 M8_UM8_4_PT5_Xo3_7(M8_UM8_4_PT5_line3, M8_UM8_4_PT5_line4, M8_UM8_4_PT5_line7);
nor2 M8_UM8_4_PT5_Xo3_8(M8_UM8_4_PT5_line5, M8_UM8_4_PT5_line6, M8_UM8_4_PT5_line8);
nand2 M8_UM8_4_PT5_Xo3_9(M8_UM8_4_PT5_line7, M8_UM8_4_PT5_line8, M8_UM8_4_line5);
inv M8_UM8_4_PT6_Xo0(M8_UM8_4_line3, M8_UM8_4_PT6_NotA);
inv M8_UM8_4_PT6_Xo1(M8_UM8_4_line4, M8_UM8_4_PT6_NotB);
nand2 M8_UM8_4_PT6_Xo2(M8_UM8_4_PT6_NotA, M8_UM8_4_line4, M8_UM8_4_PT6_line2);
nand2 M8_UM8_4_PT6_Xo3(M8_UM8_4_PT6_NotB, M8_UM8_4_line3, M8_UM8_4_PT6_line3);
nand2 M8_UM8_4_PT6_Xo4(M8_UM8_4_PT6_line2, M8_UM8_4_PT6_line3, M8_UM8_4_line6);
inv M8_UM8_4_PT7_Xo0(M8_UM8_4_line5, M8_UM8_4_PT7_NotA);
inv M8_UM8_4_PT7_Xo1(M8_UM8_4_line6, M8_UM8_4_PT7_NotB);
nand2 M8_UM8_4_PT7_Xo2(M8_UM8_4_PT7_NotA, M8_UM8_4_line6, M8_UM8_4_PT7_line2);
nand2 M8_UM8_4_PT7_Xo3(M8_UM8_4_PT7_NotB, M8_UM8_4_line5, M8_UM8_4_PT7_line3);
nand2 M8_UM8_4_PT7_Xo4(M8_UM8_4_PT7_line2, M8_UM8_4_PT7_line3, M8_ParR);
inv M8_UM8_5_PT0_Xo0(in2067, M8_UM8_5_PT0_NotA);
inv M8_UM8_5_PT0_Xo1(in2072, M8_UM8_5_PT0_NotB);
nand2 M8_UM8_5_PT0_Xo2(M8_UM8_5_PT0_NotA, in2072, M8_UM8_5_PT0_line2);
nand2 M8_UM8_5_PT0_Xo3(M8_UM8_5_PT0_NotB, in2067, M8_UM8_5_PT0_line3);
nand2 M8_UM8_5_PT0_Xo4(M8_UM8_5_PT0_line2, M8_UM8_5_PT0_line3, M8_UM8_5_line0);
inv M8_UM8_5_PT1_Xo0(in2078, M8_UM8_5_PT1_NotA);
inv M8_UM8_5_PT1_Xo1(in2084, M8_UM8_5_PT1_NotB);
nand2 M8_UM8_5_PT1_Xo2(M8_UM8_5_PT1_NotA, in2084, M8_UM8_5_PT1_line2);
nand2 M8_UM8_5_PT1_Xo3(M8_UM8_5_PT1_NotB, in2078, M8_UM8_5_PT1_line3);
nand2 M8_UM8_5_PT1_Xo4(M8_UM8_5_PT1_line2, M8_UM8_5_PT1_line3, M8_UM8_5_line1);
inv M8_UM8_5_PT2_Xo0(in2090, M8_UM8_5_PT2_NotA);
inv M8_UM8_5_PT2_Xo1(in2678, M8_UM8_5_PT2_NotB);
nand2 M8_UM8_5_PT2_Xo2(M8_UM8_5_PT2_NotA, in2678, M8_UM8_5_PT2_line2);
nand2 M8_UM8_5_PT2_Xo3(M8_UM8_5_PT2_NotB, in2090, M8_UM8_5_PT2_line3);
nand2 M8_UM8_5_PT2_Xo4(M8_UM8_5_PT2_line2, M8_UM8_5_PT2_line3, M8_UM8_5_line2);
inv M8_UM8_5_PT3_Xo0(in2100, M8_UM8_5_PT3_NotA);
inv M8_UM8_5_PT3_Xo1(in2096, M8_UM8_5_PT3_NotB);
nand2 M8_UM8_5_PT3_Xo2(M8_UM8_5_PT3_NotA, in2096, M8_UM8_5_PT3_line2);
nand2 M8_UM8_5_PT3_Xo3(M8_UM8_5_PT3_NotB, in2100, M8_UM8_5_PT3_line3);
nand2 M8_UM8_5_PT3_Xo4(M8_UM8_5_PT3_line2, M8_UM8_5_PT3_line3, M8_UM8_5_line3);
inv M8_UM8_5_PT4_Xo0(gnd, M8_UM8_5_PT4_NotA);
inv M8_UM8_5_PT4_Xo1(gnd, M8_UM8_5_PT4_NotB);
nand2 M8_UM8_5_PT4_Xo2(M8_UM8_5_PT4_NotA, gnd, M8_UM8_5_PT4_line2);
nand2 M8_UM8_5_PT4_Xo3(M8_UM8_5_PT4_NotB, gnd, M8_UM8_5_PT4_line3);
nand2 M8_UM8_5_PT4_Xo4(M8_UM8_5_PT4_line2, M8_UM8_5_PT4_line3, M8_UM8_5_line4);
inv M8_UM8_5_PT5_Xo3_0(M8_UM8_5_line0, M8_UM8_5_PT5_NotA);
inv M8_UM8_5_PT5_Xo3_1(M8_UM8_5_line1, M8_UM8_5_PT5_NotB);
inv M8_UM8_5_PT5_Xo3_2(M8_UM8_5_line2, M8_UM8_5_PT5_NotC);
and3 M8_UM8_5_PT5_Xo3_3(M8_UM8_5_PT5_NotA, M8_UM8_5_PT5_NotB, M8_UM8_5_line2, M8_UM8_5_PT5_line3);
and3 M8_UM8_5_PT5_Xo3_4(M8_UM8_5_PT5_NotA, M8_UM8_5_line1, M8_UM8_5_PT5_NotC, M8_UM8_5_PT5_line4);
and3 M8_UM8_5_PT5_Xo3_5(M8_UM8_5_line0, M8_UM8_5_PT5_NotB, M8_UM8_5_PT5_NotC, M8_UM8_5_PT5_line5);
and3 M8_UM8_5_PT5_Xo3_6(M8_UM8_5_line0, M8_UM8_5_line1, M8_UM8_5_line2, M8_UM8_5_PT5_line6);
nor2 M8_UM8_5_PT5_Xo3_7(M8_UM8_5_PT5_line3, M8_UM8_5_PT5_line4, M8_UM8_5_PT5_line7);
nor2 M8_UM8_5_PT5_Xo3_8(M8_UM8_5_PT5_line5, M8_UM8_5_PT5_line6, M8_UM8_5_PT5_line8);
nand2 M8_UM8_5_PT5_Xo3_9(M8_UM8_5_PT5_line7, M8_UM8_5_PT5_line8, M8_UM8_5_line5);
inv M8_UM8_5_PT6_Xo0(M8_UM8_5_line3, M8_UM8_5_PT6_NotA);
inv M8_UM8_5_PT6_Xo1(M8_UM8_5_line4, M8_UM8_5_PT6_NotB);
nand2 M8_UM8_5_PT6_Xo2(M8_UM8_5_PT6_NotA, M8_UM8_5_line4, M8_UM8_5_PT6_line2);
nand2 M8_UM8_5_PT6_Xo3(M8_UM8_5_PT6_NotB, M8_UM8_5_line3, M8_UM8_5_PT6_line3);
nand2 M8_UM8_5_PT6_Xo4(M8_UM8_5_PT6_line2, M8_UM8_5_PT6_line3, M8_UM8_5_line6);
inv M8_UM8_5_PT7_Xo0(M8_UM8_5_line5, M8_UM8_5_PT7_NotA);
inv M8_UM8_5_PT7_Xo1(M8_UM8_5_line6, M8_UM8_5_PT7_NotB);
nand2 M8_UM8_5_PT7_Xo2(M8_UM8_5_PT7_NotA, M8_UM8_5_line6, M8_UM8_5_PT7_line2);
nand2 M8_UM8_5_PT7_Xo3(M8_UM8_5_PT7_NotB, M8_UM8_5_line5, M8_UM8_5_PT7_line3);
nand2 M8_UM8_5_PT7_Xo4(M8_UM8_5_PT7_line2, M8_UM8_5_PT7_line3, M8_ParS);
inv M8_UM8_6(in14, M8_NotPar0);
or2 M8_UM8_7(M8_ParA, in37, M8_line7);
or2 M8_UM8_8(M8_ParB, in37, M8_line8);
or2 M8_UM8_9(M8_ParR, M8_NotPar0, M8_line9);
and3 M8_UM8_10(M8_line8, M8_line7, M8_ParS, M8_line10);
and3 M8_UM8_11(M8_ParQ, M8_line9, CompCLAs, M8_line11);
and3 M8_UM8_12(M8_line10, M8_line11, out319, out308);
inv M8_UM8_13(out308, out225);
inv M8_UM8_14(M8_line8, out395);
inv M8_UM8_15(M8_line7, out397);
inv M8_UM8_16(M8_ParS, out227);
inv M8_UM8_17(M8_ParQ, out229);
inv M8_UM8_18(M8_line9, out401);
or2 M9_UM9_0_MMC0(Abus_1, in559, M9_UM9_0_NewAbus_9);
inv M9_UM9_0_PTMuxA_PT0_Xo0(Abus_0, M9_UM9_0_PTMuxA_PT0_NotA);
inv M9_UM9_0_PTMuxA_PT0_Xo1(Abus_1, M9_UM9_0_PTMuxA_PT0_NotB);
nand2 M9_UM9_0_PTMuxA_PT0_Xo2(M9_UM9_0_PTMuxA_PT0_NotA, Abus_1, M9_UM9_0_PTMuxA_PT0_line2);
nand2 M9_UM9_0_PTMuxA_PT0_Xo3(M9_UM9_0_PTMuxA_PT0_NotB, Abus_0, M9_UM9_0_PTMuxA_PT0_line3);
nand2 M9_UM9_0_PTMuxA_PT0_Xo4(M9_UM9_0_PTMuxA_PT0_line2, M9_UM9_0_PTMuxA_PT0_line3, M9_UM9_0_PTMuxA_line0);
inv M9_UM9_0_PTMuxA_PT1_Xo0(Abus_2, M9_UM9_0_PTMuxA_PT1_NotA);
inv M9_UM9_0_PTMuxA_PT1_Xo1(Abus_5, M9_UM9_0_PTMuxA_PT1_NotB);
nand2 M9_UM9_0_PTMuxA_PT1_Xo2(M9_UM9_0_PTMuxA_PT1_NotA, Abus_5, M9_UM9_0_PTMuxA_PT1_line2);
nand2 M9_UM9_0_PTMuxA_PT1_Xo3(M9_UM9_0_PTMuxA_PT1_NotB, Abus_2, M9_UM9_0_PTMuxA_PT1_line3);
nand2 M9_UM9_0_PTMuxA_PT1_Xo4(M9_UM9_0_PTMuxA_PT1_line2, M9_UM9_0_PTMuxA_PT1_line3, M9_UM9_0_PTMuxA_line1);
inv M9_UM9_0_PTMuxA_PT2_Xo0(Abus_6, M9_UM9_0_PTMuxA_PT2_NotA);
inv M9_UM9_0_PTMuxA_PT2_Xo1(Abus_7, M9_UM9_0_PTMuxA_PT2_NotB);
nand2 M9_UM9_0_PTMuxA_PT2_Xo2(M9_UM9_0_PTMuxA_PT2_NotA, Abus_7, M9_UM9_0_PTMuxA_PT2_line2);
nand2 M9_UM9_0_PTMuxA_PT2_Xo3(M9_UM9_0_PTMuxA_PT2_NotB, Abus_6, M9_UM9_0_PTMuxA_PT2_line3);
nand2 M9_UM9_0_PTMuxA_PT2_Xo4(M9_UM9_0_PTMuxA_PT2_line2, M9_UM9_0_PTMuxA_PT2_line3, M9_UM9_0_PTMuxA_line2);
inv M9_UM9_0_PTMuxA_PT3_Xo0(Abus_8, M9_UM9_0_PTMuxA_PT3_NotA);
inv M9_UM9_0_PTMuxA_PT3_Xo1(Abus_9, M9_UM9_0_PTMuxA_PT3_NotB);
nand2 M9_UM9_0_PTMuxA_PT3_Xo2(M9_UM9_0_PTMuxA_PT3_NotA, Abus_9, M9_UM9_0_PTMuxA_PT3_line2);
nand2 M9_UM9_0_PTMuxA_PT3_Xo3(M9_UM9_0_PTMuxA_PT3_NotB, Abus_8, M9_UM9_0_PTMuxA_PT3_line3);
nand2 M9_UM9_0_PTMuxA_PT3_Xo4(M9_UM9_0_PTMuxA_PT3_line2, M9_UM9_0_PTMuxA_PT3_line3, M9_UM9_0_PTMuxA_line3);
inv M9_UM9_0_PTMuxA_PT4_Xo0(gnd, M9_UM9_0_PTMuxA_PT4_NotA);
inv M9_UM9_0_PTMuxA_PT4_Xo1(M9_UM9_0_NewAbus_9, M9_UM9_0_PTMuxA_PT4_NotB);
nand2 M9_UM9_0_PTMuxA_PT4_Xo2(M9_UM9_0_PTMuxA_PT4_NotA, M9_UM9_0_NewAbus_9, M9_UM9_0_PTMuxA_PT4_line2);
nand2 M9_UM9_0_PTMuxA_PT4_Xo3(M9_UM9_0_PTMuxA_PT4_NotB, gnd, M9_UM9_0_PTMuxA_PT4_line3);
nand2 M9_UM9_0_PTMuxA_PT4_Xo4(M9_UM9_0_PTMuxA_PT4_line2, M9_UM9_0_PTMuxA_PT4_line3, M9_UM9_0_PTMuxA_line4);
inv M9_UM9_0_PTMuxA_PT5_Xo3_0(M9_UM9_0_PTMuxA_line0, M9_UM9_0_PTMuxA_PT5_NotA);
inv M9_UM9_0_PTMuxA_PT5_Xo3_1(M9_UM9_0_PTMuxA_line1, M9_UM9_0_PTMuxA_PT5_NotB);
inv M9_UM9_0_PTMuxA_PT5_Xo3_2(M9_UM9_0_PTMuxA_line2, M9_UM9_0_PTMuxA_PT5_NotC);
and3 M9_UM9_0_PTMuxA_PT5_Xo3_3(M9_UM9_0_PTMuxA_PT5_NotA, M9_UM9_0_PTMuxA_PT5_NotB, M9_UM9_0_PTMuxA_line2, M9_UM9_0_PTMuxA_PT5_line3);
and3 M9_UM9_0_PTMuxA_PT5_Xo3_4(M9_UM9_0_PTMuxA_PT5_NotA, M9_UM9_0_PTMuxA_line1, M9_UM9_0_PTMuxA_PT5_NotC, M9_UM9_0_PTMuxA_PT5_line4);
and3 M9_UM9_0_PTMuxA_PT5_Xo3_5(M9_UM9_0_PTMuxA_line0, M9_UM9_0_PTMuxA_PT5_NotB, M9_UM9_0_PTMuxA_PT5_NotC, M9_UM9_0_PTMuxA_PT5_line5);
and3 M9_UM9_0_PTMuxA_PT5_Xo3_6(M9_UM9_0_PTMuxA_line0, M9_UM9_0_PTMuxA_line1, M9_UM9_0_PTMuxA_line2, M9_UM9_0_PTMuxA_PT5_line6);
nor2 M9_UM9_0_PTMuxA_PT5_Xo3_7(M9_UM9_0_PTMuxA_PT5_line3, M9_UM9_0_PTMuxA_PT5_line4, M9_UM9_0_PTMuxA_PT5_line7);
nor2 M9_UM9_0_PTMuxA_PT5_Xo3_8(M9_UM9_0_PTMuxA_PT5_line5, M9_UM9_0_PTMuxA_PT5_line6, M9_UM9_0_PTMuxA_PT5_line8);
nand2 M9_UM9_0_PTMuxA_PT5_Xo3_9(M9_UM9_0_PTMuxA_PT5_line7, M9_UM9_0_PTMuxA_PT5_line8, M9_UM9_0_PTMuxA_line5);
inv M9_UM9_0_PTMuxA_PT6_Xo0(M9_UM9_0_PTMuxA_line3, M9_UM9_0_PTMuxA_PT6_NotA);
inv M9_UM9_0_PTMuxA_PT6_Xo1(M9_UM9_0_PTMuxA_line4, M9_UM9_0_PTMuxA_PT6_NotB);
nand2 M9_UM9_0_PTMuxA_PT6_Xo2(M9_UM9_0_PTMuxA_PT6_NotA, M9_UM9_0_PTMuxA_line4, M9_UM9_0_PTMuxA_PT6_line2);
nand2 M9_UM9_0_PTMuxA_PT6_Xo3(M9_UM9_0_PTMuxA_PT6_NotB, M9_UM9_0_PTMuxA_line3, M9_UM9_0_PTMuxA_PT6_line3);
nand2 M9_UM9_0_PTMuxA_PT6_Xo4(M9_UM9_0_PTMuxA_PT6_line2, M9_UM9_0_PTMuxA_PT6_line3, M9_UM9_0_PTMuxA_line6);
inv M9_UM9_0_PTMuxA_PT7_Xo0(M9_UM9_0_PTMuxA_line5, M9_UM9_0_PTMuxA_PT7_NotA);
inv M9_UM9_0_PTMuxA_PT7_Xo1(M9_UM9_0_PTMuxA_line6, M9_UM9_0_PTMuxA_PT7_NotB);
nand2 M9_UM9_0_PTMuxA_PT7_Xo2(M9_UM9_0_PTMuxA_PT7_NotA, M9_UM9_0_PTMuxA_line6, M9_UM9_0_PTMuxA_PT7_line2);
nand2 M9_UM9_0_PTMuxA_PT7_Xo3(M9_UM9_0_PTMuxA_PT7_NotB, M9_UM9_0_PTMuxA_line5, M9_UM9_0_PTMuxA_PT7_line3);
nand2 M9_UM9_0_PTMuxA_PT7_Xo4(M9_UM9_0_PTMuxA_PT7_line2, M9_UM9_0_PTMuxA_PT7_line3, M9_UM9_0_ParNewA);
inv M9_UM9_0_MMC2_Mux0(in868, M9_UM9_0_MMC2_Not_ContIn);
and2 M9_UM9_0_MMC2_Mux1(Abus_9, M9_UM9_0_MMC2_Not_ContIn, M9_UM9_0_MMC2_line1);
and2 M9_UM9_0_MMC2_Mux2(M9_UM9_0_ParNewA, in868, M9_UM9_0_MMC2_line2);
or2 M9_UM9_0_MMC2_Mux3(M9_UM9_0_MMC2_line1, M9_UM9_0_MMC2_line2, out331);
inv M9_UM9_0_MMC3_Mux0(in868, M9_UM9_0_MMC3_Not_ContIn);
and2 M9_UM9_0_MMC3_Mux1(Abus_0, M9_UM9_0_MMC3_Not_ContIn, M9_UM9_0_MMC3_line1);
and2 M9_UM9_0_MMC3_Mux2(M9_UM9_0_NewAbus_9, in868, M9_UM9_0_MMC3_line2);
or2 M9_UM9_0_MMC3_Mux3(M9_UM9_0_MMC3_line1, M9_UM9_0_MMC3_line2, out323);
inv M9_UM9_0_MMC4_Mux0(in868, M9_UM9_0_MMC4_Not_ContIn);
and2 M9_UM9_0_MMC4_Mux1(Abus_1, M9_UM9_0_MMC4_Not_ContIn, M9_UM9_0_MMC4_line1);
and2 M9_UM9_0_MMC4_Mux2(Abus_3, in868, M9_UM9_0_MMC4_line2);
or2 M9_UM9_0_MMC4_Mux3(M9_UM9_0_MMC4_line1, M9_UM9_0_MMC4_line2, out321);
inv M9_UM9_0_MMC5_Mux0(in868, M9_UM9_0_MMC5_Not_ContIn);
and2 M9_UM9_0_MMC5_Mux1(Abus_2, M9_UM9_0_MMC5_Not_ContIn, M9_UM9_0_MMC5_line1);
and2 M9_UM9_0_MMC5_Mux2(Abus_4, in868, M9_UM9_0_MMC5_line2);
or2 M9_UM9_0_MMC5_Mux3(M9_UM9_0_MMC5_line1, M9_UM9_0_MMC5_line2, out280);
inv M9_UM9_0_MMC6(M9_UM9_0_NewAbus_9, M9_UM9_0_NotNewA9);
inv M9_UM9_0_MMC7_Xo0(Abus_0, M9_UM9_0_MMC7_NotA);
inv M9_UM9_0_MMC7_Xo1(Abus_1, M9_UM9_0_MMC7_NotB);
nand2 M9_UM9_0_MMC7_Xo2(M9_UM9_0_MMC7_NotA, Abus_1, M9_UM9_0_MMC7_line2);
nand2 M9_UM9_0_MMC7_Xo3(M9_UM9_0_MMC7_NotB, Abus_0, M9_UM9_0_MMC7_line3);
nand2 M9_UM9_0_MMC7_Xo4(M9_UM9_0_MMC7_line2, M9_UM9_0_MMC7_line3, M9_UM9_0_line7);
inv M9_UM9_0_MMC8_Xo0(M9_UM9_0_line7, M9_UM9_0_MMC8_NotA);
inv M9_UM9_0_MMC8_Xo1(M9_UM9_0_NotNewA9, M9_UM9_0_MMC8_NotB);
nand2 M9_UM9_0_MMC8_Xo2(M9_UM9_0_MMC8_NotA, M9_UM9_0_NotNewA9, M9_UM9_0_MMC8_line2);
nand2 M9_UM9_0_MMC8_Xo3(M9_UM9_0_MMC8_NotB, M9_UM9_0_line7, M9_UM9_0_MMC8_line3);
nand2 M9_UM9_0_MMC8_Xo4(M9_UM9_0_MMC8_line2, M9_UM9_0_MMC8_line3, M9_UM9_0_line8);
inv M9_UM9_0_MMC9_Xo0(M9_UM9_0_line8, M9_UM9_0_MMC9_NotA);
inv M9_UM9_0_MMC9_Xo1(Abus_9, M9_UM9_0_MMC9_NotB);
nand2 M9_UM9_0_MMC9_Xo2(M9_UM9_0_MMC9_NotA, Abus_9, M9_UM9_0_MMC9_line2);
nand2 M9_UM9_0_MMC9_Xo3(M9_UM9_0_MMC9_NotB, M9_UM9_0_line8, M9_UM9_0_MMC9_line3);
nand2 M9_UM9_0_MMC9_Xo4(M9_UM9_0_MMC9_line2, M9_UM9_0_MMC9_line3, M9_UM9_0_line9);
inv M9_UM9_0_MMC10_Mux0(in860, M9_UM9_0_MMC10_Not_ContIn);
and2 M9_UM9_0_MMC10_Mux1(M9_UM9_0_line9, M9_UM9_0_MMC10_Not_ContIn, M9_UM9_0_MMC10_line1);
and2 M9_UM9_0_MMC10_Mux2(Abus_9, in860, M9_UM9_0_MMC10_line2);
or2 M9_UM9_0_MMC10_Mux3(M9_UM9_0_MMC10_line1, M9_UM9_0_MMC10_line2, out145);
inv M9_UM9_0_MMC11_Mux0(in860, M9_UM9_0_MMC11_Not_ContIn);
and2 M9_UM9_0_MMC11_Mux1(M9_UM9_0_NewAbus_9, M9_UM9_0_MMC11_Not_ContIn, M9_UM9_0_MMC11_line1);
and2 M9_UM9_0_MMC11_Mux2(Abus_1, in860, M9_UM9_0_MMC11_line2);
or2 M9_UM9_0_MMC11_Mux3(M9_UM9_0_MMC11_line1, M9_UM9_0_MMC11_line2, out148);
inv M9_UM9_0_MMC12_Mux0(in860, M9_UM9_0_MMC12_Not_ContIn);
and2 M9_UM9_0_MMC12_Mux1(vdd, M9_UM9_0_MMC12_Not_ContIn, M9_UM9_0_MMC12_line1);
and2 M9_UM9_0_MMC12_Mux2(Abus_0, in860, M9_UM9_0_MMC12_line2);
or2 M9_UM9_0_MMC12_Mux3(M9_UM9_0_MMC12_line1, M9_UM9_0_MMC12_line2, out153);
buffer M9_UM9_1_MBC0(Abus_8, out290);
buffer M9_UM9_1_MBC1(Abus_7, out305);
buffer M9_UM9_1_MBC2(Abus_6, out288);
buffer M9_UM9_1_MBC3(Abus_5, out303);
buffer M9_UM9_1_MBC4(Abus_4, out286);
buffer M9_UM9_1_MBC5(Abus_3, out301);
buffer M9_UM9_1_MBC6(Abus_2, out299);
inv M9_UM9_1_MBC7(Abus_5, out166);
inv M9_UM9_1_MBC8(Abus_4, out168);
inv M9_UM9_1_MBC9(Abus_3, out171);
inv M9_UM9_1_MBC10(Bbus_6, out162);
inv M9_UM9_1_MBC11(Bbus_5, out160);
inv M9_UM9_1_MBC12(Bbus_4, out164);
buffer M9_UM9_2_MRC0(in452, out335);
buffer M9_UM9_2_MRC1(in452, out350);
buffer M9_UM9_2_MRC2(in452, out391);
buffer M9_UM9_2_MRC3(in452, out409);
buffer M9_UM9_2_MRC4(in2066, out337);
buffer M9_UM9_2_MRC5(in2066, out384);
buffer M9_UM9_2_MRC6(in2066, out411);
buffer M9_UM9_2_MRC7(in1083, out367);
buffer M9_UM9_2_MRC8(in1083, out369);
and2 M9_UM9_2_MRC9(in452, in94, out173);
inv M9_UM9_2_MRC10(in2100, M9_UM9_2_NotPTIns10);
inv M9_UM9_2_MRC11(in2096, M9_UM9_2_NotPTIns11);
nand2 M9_UM9_2_MRC12_Xo1_0(Bbus_9, M9_UM9_2_NotPTIns10, M9_UM9_2_MRC12_NotAB);
and2 M9_UM9_2_MRC12_Xo1_1(Bbus_9, M9_UM9_2_MRC12_NotAB, M9_UM9_2_MRC12_line1);
and2 M9_UM9_2_MRC12_Xo1_2(M9_UM9_2_MRC12_NotAB, M9_UM9_2_NotPTIns10, M9_UM9_2_MRC12_line2);
or2 M9_UM9_2_MRC12_Xo1_3(M9_UM9_2_MRC12_line1, M9_UM9_2_MRC12_line2, M9_UM9_2_line12);
nand2 M9_UM9_2_MRC13_Xo1_0(Bbus_7, M9_UM9_2_NotPTIns11, M9_UM9_2_MRC13_NotAB);
and2 M9_UM9_2_MRC13_Xo1_1(Bbus_7, M9_UM9_2_MRC13_NotAB, M9_UM9_2_MRC13_line1);
and2 M9_UM9_2_MRC13_Xo1_2(M9_UM9_2_MRC13_NotAB, M9_UM9_2_NotPTIns11, M9_UM9_2_MRC13_line2);
or2 M9_UM9_2_MRC13_Xo1_3(M9_UM9_2_MRC13_line1, M9_UM9_2_MRC13_line2, M9_UM9_2_line13);
inv M9_UM9_2_MRC14_RIV0(M9_UM9_2_line12, M9_UM9_2_MRC14_NotA);
and2 M9_UM9_2_MRC14_RIV1(M9_UM9_2_line12, M9_UM9_2_MRC14_NotA, M9_UM9_2_MRC14_line1);
or2 M9_UM9_2_MRC14_RIV2(M9_UM9_2_MRC14_line1, M9_UM9_2_MRC14_NotA, M9_UM9_2_line14);
inv M9_UM9_2_MRC15_RIV0(M9_UM9_2_line13, M9_UM9_2_MRC15_NotA);
and2 M9_UM9_2_MRC15_RIV1(M9_UM9_2_line13, M9_UM9_2_MRC15_NotA, M9_UM9_2_MRC15_line1);
or2 M9_UM9_2_MRC15_RIV2(M9_UM9_2_MRC15_line1, M9_UM9_2_MRC15_NotA, M9_UM9_2_line15);
nand2 M9_UM9_2_MRC16(M9_UM9_2_line14, M9_UM9_2_line15, out156);
and2 M9_UM9_2_MRC17(in7, in661, M9_UM9_2_line17);
inv M9_UM9_2_MRC18(M9_UM9_2_line17, out223);
and2 M9_UM9_2_MRC19(in2106, M9_UM9_2_line17, M9_UM9_2_line19);
inv M9_UM9_2_MRC20(M9_UM9_2_line19, out217);
nand2 M9_UM9_2_MRC21(in567, M9_UM9_2_line17, out234);
and3 M9_UM9_2_MRC22(in2, in15, in661, M9_UM9_2_line22);
inv M9_UM9_2_MRC23(M9_UM9_2_line22, out259);
and4 M9_UM9_2_MRC24(in661, in483, in36, out319, M9_UM9_2_line24);
inv M9_UM9_2_MRC25(M9_UM9_2_line24, out176);
and2 M9_UM9_2_MRC26(in1, in3, M9_UM9_2_line26);
inv M9_UM9_2_MRC27(M9_UM9_2_line26, M9_UM9_2_line27);
and4 M9_UM9_2_MRC28(in661, in483, out319, M9_UM9_2_line27, M9_UM9_2_line28);
inv M9_UM9_2_MRC29(M9_UM9_2_line28, out188);
and4 M9_UM9_2_MRC30(in2072, in2078, in2084, in2090, M9_UM9_2_line30);
inv M9_UM9_2_MRC31(M9_UM9_2_line30, out158);

assign out295 = out331;
assign out282 = out323;
assign out284 = out321;
assign out297 = out280;
assign out169 = in169;
assign out174 = in174;
assign out177 = in177;
assign out178 = in178;
assign out179 = in179;
assign out180 = in180;
assign out181 = in181;
assign out182 = in182;
assign out183 = in183;
assign out184 = in184;
assign out185 = in185;
assign out186 = in186;
assign out189 = in189;
assign out190 = in190;
assign out191 = in191;
assign out192 = in192;
assign out193 = in193;
assign out194 = in194;
assign out195 = in195;
assign out196 = in196;
assign out197 = in197;
assign out198 = in198;
assign out199 = in199;
assign out200 = in200;
assign out201 = in201;
assign out202 = in202;
assign out203 = in203;
assign out204 = in204;
assign out205 = in205;
assign out206 = in206;
assign out207 = in207;
assign out208 = in208;
assign out209 = in209;
assign out210 = in210;
assign out211 = in211;
assign out212 = in212;
assign out213 = in213;
assign out214 = in214;
assign out215 = in215;
assign out239 = in239;
assign out240 = in240;
assign out241 = in241;
assign out242 = in242;
assign out243 = in243;
assign out244 = in244;
assign out245 = in245;
assign out246 = in246;
assign out247 = in247;
assign out248 = in248;
assign out249 = in249;
assign out250 = in250;
assign out251 = in251;
assign out252 = in252;
assign out253 = in253;
assign out254 = in254;
assign out255 = in255;
assign out256 = in256;
assign out257 = in257;
assign out262 = in262;
assign out263 = in263;
assign out264 = in264;
assign out265 = in265;
assign out266 = in266;
assign out267 = in267;
assign out268 = in268;
assign out269 = in269;
assign out270 = in270;
assign out271 = in271;
assign out272 = in272;
assign out273 = in273;
assign out274 = in274;
assign out275 = in275;
assign out276 = in276;
assign out277 = in277;
assign out278 = in278;
assign out279 = in279;
assign vdd = 1'b1;
assign gnd = 1'b0;

endmodule
