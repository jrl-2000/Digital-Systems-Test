module c1908(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G1884,G1885,G1886,G1887,
  G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G19,
  G1900,G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G2,G20,G21,G22,G23,G24,
  G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G4,G5,G6,G7,G8,G9);
  
input G1;
input G2;
input G3;
input G4;
input G5;
input G6;
input G7;
input G8;
input G9;
input G10;
input G11;
input G12;
input G13;
input G14;
input G15;
input G16;
input G17;
input G18;
input G19;
input G20;
input G21;
input G22;
input G23;
input G24;
input G25;
input G26;
input G27;
input G28;
input G29;
input G30;
input G31;
input G32;
input G33;

output G1884;
output G1885;
output G1886;
output G1887;
output G1888;
output G1889;
output G1890;
output G1891;
output G1892;
output G1893;
output G1894;
output G1895;
output G1896;
output G1897;
output G1898;
output G1899;
output G1900;
output G1901;
output G1902;
output G1903;
output G1904;
output G1905;
output G1906;
output G1907;
output G1908;

  wire G112,G116,G119,G123,G128,G131,G134,G138,G142,G147,G151,G154,G157,G161,
    G165,G169,G173,G174,G175,G178,G179,G182,G185,G188,G191,G194,G197,G198,G199,
    G202,G205,G212,G219,G222,G225,G228,G235,G238,G241,G248,G253,G260,G265,G268,
    G271,G274,G277,G280,G283,G286,G289,G292,G295,G298,G301,G304,G307,G310,G313,
    G314,G315,G316,G317,G318,G319,G320,G321,G322,G323,G324,G325,G326,G327,G328,
    G329,G330,G331,G332,G333,G334,G335,G338,G341,G344,G347,G350,G353,G356,G359,
    G362,G365,G368,G371,G374,G377,G380,G381,G382,G387,G391,G395,G398,G401,G404,
    G407,G410,G413,G416,G419,G422,G425,G428,G431,G434,G437,G440,G443,G446,G449,
    G452,G455,G458,G461,G464,G467,G470,G473,G476,G479,G482,G485,G488,G491,G494,
    G497,G500,G503,G506,G509,G512,G515,G518,G521,G524,G527,G530,G533,G534,G535,
    G536,G537,G538,G539,G540,G541,G542,G543,G544,G545,G546,G550,G554,G557,G560,
    G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G573,G582,G585,G586,G589,
    G590,G593,G594,G597,G598,G601,G602,G605,G606,G609,G612,G615,G616,G619,G620,
    G623,G624,G627,G628,G631,G632,G635,G636,G637,G638,G639,G640,G641,G644,G645,
    G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G660,G663,G666,G669,G672,
    G675,G678,G681,G684,G687,G690,G693,G696,G699,G700,G701,G702,G703,G704,G705,
    G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
    G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G734,G735,G738,G755,
    G772,G773,G774,G775,G776,G777,G778,G779,G780,G781,G782,G783,G784,G785,G786,
    G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G802,G805,
    G806,G807,G808,G809,G810,G813,G816,G819,G822,G825,G828,G831,G834,G835,G836,
    G837,G838,G839,G840,G841,G842,G843,G844,G845,G848,G849,G850,G851,G854,G855,
    G856,G857,G858,G859,G860,G861,G864,G867,G870,G873,G876,G879,G882,G885,G888,
    G891,G894,G895,G896,G897,G898,G901,G904,G905,G906,G907,G908,G909,G910,G911,
    G914,G917,G918,G919,G920,G921,G924,G925,G926,G927,G928,G929,G930,G931,G932,
    G933,G934,G935,G936,G937,G938,G939,G940,G941,G942,G943,G944,G945,G946,G947,
    G948,G951,G952,G953,G956,G959,G962,G963,G964,G965,G966,G967,G968,G969,G970,
    G971,G972,G973,G974,G975,G976,G977,G980,G981,G984,G987,G988,G989,G993,G994,
    G995,G996,G997,G998,G999,G1000,G1003,G1006,G1009,G1012,G1015,G1019,G1022,
    G1023,G1024,G1025,G1028,G1031,G1034,G1035,G1036,G1037,G1038,G1041,G1044,
    G1047,G1050,G1053,G1056,G1059,G1062,G1065,G1066,G1067,G1068,G1069,G1072,
    G1075,G1078,G1081,G1084,G1087,G1090,G1091,G1092,G1093,G1094,G1095,G1096,
    G1097,G1098,G1099,G1100,G1103,G1104,G1107,G1110,G1111,G1112,G1113,G1114,
    G1115,G1116,G1117,G1118,G1121,G1124,G1125,G1126,G1129,G1130,G1131,G1132,
    G1135,G1138,G1139,G1140,G1143,G1144,G1145,G1148,G1151,G1152,G1153,G1154,
    G1155,G1156,G1157,G1158,G1159,G1160,G1163,G1166,G1167,G1168,G1169,G1170,
    G1171,G1174,G1175,G1176,G1177,G1178,G1181,G1182,G1185,G1186,G1187,G1188,
    G1189,G1192,G1195,G1198,G1199,G1200,G1201,G1202,G1203,G1204,G1205,G1208,
    G1209,G1212,G1215,G1216,G1217,G1218,G1219,G1220,G1221,G1222,G1225,G1226,
    G1227,G1230,G1233,G1236,G1239,G1240,G1243,G1244,G1245,G1246,G1247,G1250,
    G1251,G1252,G1253,G1256,G1259,G1260,G1261,G1262,G1263,G1264,G1265,G1266,
    G1267,G1268,G1269,G1270,G1273,G1276,G1279,G1280,G1281,G1282,G1283,G1284,
    G1287,G1290,G1293,G1296,G1299,G1302,G1305,G1308,G1309,G1310,G1311,G1312,
    G1313,G1316,G1317,G1320,G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,
    G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
    G1341,G1342,G1343,G1344,G1347,G1350,G1353,G1354,G1355,G1356,G1357,G1358,
    G1359,G1362,G1363,G1366,G1369,G1370,G1371,G1374,G1375,G1378,G1381,G1382,
    G1383,G1386,G1389,G1392,G1395,G1410,G1420,G1434,G1439,G1442,G1445,G1448,
    G1451,G1454,G1457,G1458,G1459,G1460,G1461,G1462,G1463,G1464,G1465,G1466,
    G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1479,G1480,
    G1483,G1484,G1487,G1488,G1489,G1490,G1493,G1496,G1499,G1502,G1505,G1508,
    G1511,G1522,G1538,G1549,G1563,G1576,G1584,G1598,G1607,G1608,G1609,G1624,
    G1625,G1642,G1645,G1648,G1651,G1654,G1657,G1660,G1663,G1666,G1669,G1672,
    G1675,G1678,G1681,G1684,G1687,G1690,G1693,G1696,G1699,G1702,G1705,G1708,
    G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1722,G1725,G1728,
    G1731,G1734,G1737,G1740,G1743,G1746,G1747,G1748,G1749,G1750,G1751,G1752,
    G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,G1761,G1762,G1763,G1764,
    G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,
    G1777,G1778,G1779,G1780,G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,
    G1791,G1794,G1795,G1796,G1797,G1798,G1799,G1800,G1801,G1802,G1803,G1806,
    G1809,G1810,G1817,G1818,G1819,G1820,G1821,G1822,G1825,G1828,G1831,G1834,
    G1837,G1838,G1839,G1842,G1845,G1848,G1849,G1850,G1851,G1852,G1853,G1854,
    G1855,G1856,G1857,G1858,G1859,G1860,G1861,G1862,G1863,G1864,G1865,G1866,
    G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1880,
    G1881,G1882,G1883;

  not NOT_0(G112,G1);
  not NOT_1(G116,G2);
  not NOT_2(G119,G3);
  not NOT_3(G123,G4);
  not NOT_4(G128,G5);
  not NOT_5(G131,G6);
  not NOT_6(G134,G7);
  not NOT_7(G138,G8);
  not NOT_8(G142,G9);
  not NOT_9(G147,G10);
  not NOT_10(G151,G11);
  not NOT_11(G154,G12);
  not NOT_12(G157,G13);
  not NOT_13(G161,G14);
  not NOT_14(G165,G15);
  not NOT_15(G169,G16);
  nand NAND2_0(G173,G21,G29);
  nand NAND2_1(G174,G22,G30);
  not NOT_16(G175,G24);
  not NOT_17(G178,G24);
  not NOT_18(G179,G23);
  not NOT_19(G182,G23);
  not NOT_20(G185,G25);
  not NOT_21(G188,G26);
  not NOT_22(G191,G27);
  not NOT_23(G194,G28);
  not NOT_24(G197,G33);
  not NOT_25(G198,G33);
  not NOT_26(G199,G29);
  not NOT_27(G202,G30);
  not NOT_28(G205,G31);
  not NOT_29(G212,G31);
  not NOT_30(G219,G31);
  not NOT_31(G222,G31);
  not NOT_32(G225,G32);
  not NOT_33(G228,G32);
  not NOT_34(G235,G32);
  not NOT_35(G238,G33);
  not NOT_36(G241,G33);
  not NOT_37(G248,G33);
  not NOT_38(G253,G33);
  not NOT_39(G260,G33);
  not NOT_40(G265,G1);
  not NOT_41(G268,G2);
  not NOT_42(G271,G3);
  not NOT_43(G274,G4);
  not NOT_44(G277,G5);
  not NOT_45(G280,G6);
  not NOT_46(G283,G7);
  not NOT_47(G286,G8);
  not NOT_48(G289,G9);
  not NOT_49(G292,G10);
  not NOT_50(G295,G11);
  not NOT_51(G298,G12);
  not NOT_52(G301,G13);
  not NOT_53(G304,G14);
  not NOT_54(G307,G15);
  not NOT_55(G310,G16);
  not NOT_56(G313,G265);
  not NOT_57(G314,G268);
  not NOT_58(G315,G271);
  not NOT_59(G316,G274);
  not NOT_60(G317,G277);
  not NOT_61(G318,G280);
  not NOT_62(G319,G283);
  not NOT_63(G320,G286);
  not NOT_64(G321,G289);
  not NOT_65(G322,G292);
  not NOT_66(G323,G295);
  not NOT_67(G324,G298);
  not NOT_68(G325,G301);
  not NOT_69(G326,G304);
  not NOT_70(G327,G307);
  not NOT_71(G328,G310);
  nand NAND2_2(G329,G228,G253);
  nand NAND2_3(G330,G228,G253);
  nand NAND2_4(G331,G228,G253);
  nand NAND2_5(G332,G228,G253);
  nand NAND2_6(G333,G228,G253);
  nand NAND2_7(G334,G228,G253);
  not NOT_72(G335,G112);
  not NOT_73(G338,G116);
  not NOT_74(G341,G128);
  not NOT_75(G344,G131);
  not NOT_76(G347,G147);
  not NOT_77(G350,G165);
  and AND2_0(G353,G21,G241);
  not NOT_78(G356,G142);
  not NOT_79(G359,G151);
  not NOT_80(G362,G154);
  and AND2_1(G365,G22,G241);
  not NOT_81(G368,G161);
  and AND3_0(G371,G17,G175,G241);
  not NOT_82(G374,G169);
  not NOT_83(G377,G161);
  nand NAND2_8(G380,G248,G199);
  nand NAND2_9(G381,G248,G202);
  nand NAND2_10(G382,G182,G24);
  nand NAND2_11(G387,G182,G222);
  nand NAND2_12(G391,G178,G222);
  not NOT_84(G395,G123);
  not NOT_85(G398,G138);
  not NOT_86(G401,G142);
  not NOT_87(G404,G161);
  not NOT_88(G407,G112);
  not NOT_89(G410,G112);
  not NOT_90(G413,G116);
  not NOT_91(G416,G151);
  not NOT_92(G419,G119);
  and AND3_1(G422,G19,G179,G241);
  not NOT_93(G425,G154);
  not NOT_94(G428,G123);
  not NOT_95(G431,G157);
  and AND3_2(G434,G20,G179,G241);
  not NOT_96(G437,G185);
  not NOT_97(G440,G185);
  not NOT_98(G443,G188);
  not NOT_99(G446,G188);
  not NOT_100(G449,G191);
  not NOT_101(G452,G191);
  not NOT_102(G455,G194);
  not NOT_103(G458,G194);
  and AND2_2(G461,G173,G238);
  and AND2_3(G464,G174,G238);
  not NOT_104(G467,G119);
  not NOT_105(G470,G119);
  not NOT_106(G473,G134);
  not NOT_107(G476,G134);
  not NOT_108(G479,G169);
  not NOT_109(G482,G169);
  not NOT_110(G485,G157);
  not NOT_111(G488,G157);
  not NOT_112(G491,G123);
  not NOT_113(G494,G123);
  not NOT_114(G497,G128);
  not NOT_115(G500,G138);
  and AND3_3(G503,G18,G175,G241);
  not NOT_116(G506,G165);
  not NOT_117(G509,G142);
  not NOT_118(G512,G142);
  not NOT_119(G515,G131);
  not NOT_120(G518,G138);
  not NOT_121(G521,G147);
  not NOT_122(G524,G165);
  not NOT_123(G527,G134);
  not NOT_124(G530,G147);
  not NOT_125(G533,G461);
  not NOT_126(G534,G464);
  not NOT_127(G535,G395);
  not NOT_128(G536,G398);
  not NOT_129(G537,G401);
  not NOT_130(G538,G404);
  not NOT_131(G539,G410);
  not NOT_132(G540,G422);
  not NOT_133(G541,G428);
  not NOT_134(G542,G431);
  not NOT_135(G543,G434);
  and AND2_4(G544,G17,G391);
  and AND2_5(G545,G19,G387);
  nand NAND2_13(G546,G18,G391);
  nand NAND2_14(G550,G20,G387);
  nand NAND2_15(G554,G17,G391);
  nand NAND2_16(G557,G19,G387);
  not NOT_136(G560,G440);
  not NOT_137(G561,G437);
  not NOT_138(G562,G446);
  not NOT_139(G563,G443);
  not NOT_140(G564,G452);
  not NOT_141(G565,G449);
  not NOT_142(G566,G458);
  not NOT_143(G567,G455);
  nand NAND4_0(G568,G199,G219,G248,G382);
  nand NAND4_1(G569,G202,G219,G248,G382);
  nand NAND3_0(G570,G225,G260,G382);
  and AND3_4(G573,G225,G260,G382);
  not NOT_144(G582,G335);
  not NOT_145(G585,G467);
  not NOT_146(G586,G335);
  not NOT_147(G589,G470);
  not NOT_148(G590,G341);
  not NOT_149(G593,G473);
  not NOT_150(G594,G341);
  not NOT_151(G597,G476);
  not NOT_152(G598,G347);
  not NOT_153(G601,G479);
  not NOT_154(G602,G347);
  not NOT_155(G605,G482);
  not NOT_156(G606,G353);
  not NOT_157(G609,G353);
  not NOT_158(G612,G359);
  not NOT_159(G615,G485);
  not NOT_160(G616,G359);
  not NOT_161(G619,G488);
  not NOT_162(G620,G365);
  not NOT_163(G623,G491);
  not NOT_164(G624,G365);
  not NOT_165(G627,G494);
  not NOT_166(G628,G371);
  not NOT_167(G631,G407);
  not NOT_168(G632,G371);
  not NOT_169(G635,G497);
  not NOT_170(G636,G500);
  not NOT_171(G637,G413);
  not NOT_172(G638,G503);
  not NOT_173(G639,G506);
  not NOT_174(G640,G416);
  not NOT_175(G641,G374);
  not NOT_176(G644,G509);
  not NOT_177(G645,G374);
  not NOT_178(G648,G512);
  not NOT_179(G649,G515);
  not NOT_180(G650,G518);
  not NOT_181(G651,G419);
  not NOT_182(G652,G521);
  not NOT_183(G653,G524);
  not NOT_184(G654,G425);
  not NOT_185(G655,G527);
  not NOT_186(G656,G530);
  not NOT_187(G657,G338);
  not NOT_188(G660,G338);
  not NOT_189(G663,G344);
  not NOT_190(G666,G344);
  not NOT_191(G669,G350);
  not NOT_192(G672,G350);
  not NOT_193(G675,G356);
  not NOT_194(G678,G356);
  not NOT_195(G681,G362);
  not NOT_196(G684,G362);
  not NOT_197(G687,G368);
  not NOT_198(G690,G368);
  not NOT_199(G693,G377);
  not NOT_200(G696,G377);
  nand NAND2_17(G699,G398,G535);
  nand NAND2_18(G700,G395,G536);
  nand NAND2_19(G701,G404,G537);
  nand NAND2_20(G702,G401,G538);
  nand NAND2_21(G703,G434,G542);
  nand NAND2_22(G704,G431,G543);
  nand NAND2_23(G705,G500,G635);
  nand NAND2_24(G706,G497,G636);
  nand NAND2_25(G707,G506,G638);
  nand NAND2_26(G708,G503,G639);
  nand NAND2_27(G709,G518,G649);
  nand NAND2_28(G710,G515,G650);
  nand NAND2_29(G711,G524,G652);
  nand NAND2_30(G712,G521,G653);
  nand NAND2_31(G713,G530,G655);
  nand NAND2_32(G714,G527,G656);
  not NOT_201(G715,G586);
  not NOT_202(G716,G582);
  nand NAND2_33(G717,G699,G700);
  not NOT_203(G718,G590);
  not NOT_204(G719,G594);
  not NOT_205(G720,G602);
  not NOT_206(G721,G598);
  not NOT_207(G722,G609);
  not NOT_208(G723,G616);
  not NOT_209(G724,G624);
  nand NAND2_34(G725,G701,G702);
  not NOT_210(G726,G632);
  nand NAND2_35(G727,G632,G539);
  not NOT_211(G728,G645);
  nand NAND2_36(G729,G703,G704);
  not NOT_212(G730,G546);
  not NOT_213(G731,G546);
  not NOT_214(G734,G550);
  not NOT_215(G735,G550);
  nand NAND2_37(G738,G568,G570);
  nand NAND2_38(G755,G569,G570);
  not NOT_216(G772,G657);
  nand NAND2_39(G773,G657,G585);
  not NOT_217(G774,G660);
  nand NAND2_40(G775,G660,G589);
  not NOT_218(G776,G663);
  nand NAND2_41(G777,G663,G593);
  not NOT_219(G778,G666);
  nand NAND2_42(G779,G666,G597);
  not NOT_220(G780,G669);
  nand NAND2_43(G781,G669,G601);
  not NOT_221(G782,G672);
  nand NAND2_44(G783,G672,G605);
  not NOT_222(G784,G675);
  not NOT_223(G785,G606);
  not NOT_224(G786,G678);
  not NOT_225(G787,G681);
  nand NAND2_45(G788,G681,G615);
  not NOT_226(G789,G612);
  not NOT_227(G790,G684);
  nand NAND2_46(G791,G684,G619);
  not NOT_228(G792,G687);
  nand NAND2_47(G793,G687,G623);
  not NOT_229(G794,G620);
  not NOT_230(G795,G690);
  nand NAND2_48(G796,G690,G627);
  not NOT_231(G797,G628);
  nand NAND2_49(G798,G628,G631);
  nand NAND2_50(G799,G705,G706);
  nand NAND2_51(G802,G707,G708);
  not NOT_232(G805,G693);
  nand NAND2_52(G806,G693,G644);
  not NOT_233(G807,G641);
  not NOT_234(G808,G696);
  nand NAND2_53(G809,G696,G648);
  nand NAND2_54(G810,G709,G710);
  nand NAND2_55(G813,G711,G712);
  nand NAND2_56(G816,G713,G714);
  not NOT_235(G819,G554);
  not NOT_236(G822,G554);
  not NOT_237(G825,G557);
  not NOT_238(G828,G557);
  not NOT_239(G831,G717);
  nand NAND2_57(G834,G410,G726);
  nand NAND2_58(G835,G467,G772);
  nand NAND2_59(G836,G470,G774);
  nand NAND2_60(G837,G473,G776);
  nand NAND2_61(G838,G476,G778);
  nand NAND2_62(G839,G479,G780);
  nand NAND2_63(G840,G482,G782);
  nand NAND2_64(G841,G485,G787);
  nand NAND2_65(G842,G488,G790);
  nand NAND2_66(G843,G491,G792);
  nand NAND2_67(G844,G494,G795);
  not NOT_240(G845,G725);
  nand NAND2_68(G848,G407,G797);
  nand NAND2_69(G849,G509,G805);
  nand NAND2_70(G850,G512,G808);
  not NOT_241(G851,G729);
  nand NAND2_71(G854,G834,G727);
  nand NAND2_72(G855,G816,G541);
  not NOT_242(G856,G816);
  not NOT_243(G857,G822);
  not NOT_244(G858,G819);
  not NOT_245(G859,G828);
  not NOT_246(G860,G825);
  nand NAND2_73(G861,G835,G773);
  nand NAND2_74(G864,G836,G775);
  nand NAND2_75(G867,G837,G777);
  nand NAND2_76(G870,G838,G779);
  nand NAND2_77(G873,G839,G781);
  nand NAND2_78(G876,G840,G783);
  nand NAND2_79(G879,G841,G788);
  nand NAND2_80(G882,G842,G791);
  nand NAND2_81(G885,G843,G793);
  nand NAND2_82(G888,G844,G796);
  nand NAND2_83(G891,G848,G798);
  not NOT_247(G894,G799);
  nand NAND2_84(G895,G799,G637);
  not NOT_248(G896,G802);
  nand NAND2_85(G897,G802,G640);
  nand NAND2_86(G898,G849,G806);
  nand NAND2_87(G901,G850,G809);
  not NOT_249(G904,G810);
  nand NAND2_88(G905,G810,G651);
  not NOT_250(G906,G813);
  nand NAND2_89(G907,G813,G654);
  not NOT_251(G908,G845);
  nand NAND2_90(G909,G428,G856);
  not NOT_252(G910,G851);
  not NOT_253(G911,G831);
  not NOT_254(G914,G831);
  nand NAND2_91(G917,G413,G894);
  nand NAND2_92(G918,G416,G896);
  nand NAND2_93(G919,G419,G904);
  nand NAND2_94(G920,G425,G906);
  not NOT_255(G921,G854);
  nand NAND2_95(G924,G864,G715);
  not NOT_256(G925,G864);
  nand NAND2_96(G926,G861,G716);
  not NOT_257(G927,G861);
  nand NAND2_97(G928,G867,G718);
  not NOT_258(G929,G867);
  nand NAND2_98(G930,G870,G719);
  not NOT_259(G931,G870);
  nand NAND2_99(G932,G876,G720);
  not NOT_260(G933,G876);
  nand NAND2_100(G934,G873,G721);
  not NOT_261(G935,G873);
  nand NAND2_101(G936,G882,G723);
  not NOT_262(G937,G882);
  nand NAND2_102(G938,G888,G724);
  not NOT_263(G939,G888);
  not NOT_264(G940,G891);
  nand NAND2_103(G941,G901,G728);
  not NOT_265(G942,G901);
  nand NAND2_104(G943,G855,G909);
  not NOT_266(G944,G879);
  nand NAND2_105(G945,G879,G789);
  not NOT_267(G946,G885);
  nand NAND2_106(G947,G885,G794);
  nand NAND2_107(G948,G895,G917);
  not NOT_268(G951,G898);
  nand NAND2_108(G952,G898,G807);
  nand NAND2_109(G953,G897,G918);
  nand NAND2_110(G956,G907,G920);
  nand NAND2_111(G959,G905,G919);
  nand NAND2_112(G962,G586,G925);
  nand NAND2_113(G963,G582,G927);
  nand NAND2_114(G964,G590,G929);
  not NOT_269(G965,G914);
  not NOT_270(G966,G911);
  nand NAND2_115(G967,G594,G931);
  nand NAND2_116(G968,G602,G933);
  nand NAND2_117(G969,G598,G935);
  nand NAND2_118(G970,G616,G937);
  nand NAND2_119(G971,G624,G939);
  nand NAND2_120(G972,G645,G942);
  not NOT_271(G973,G921);
  nand NAND2_121(G974,G612,G944);
  nand NAND2_122(G975,G620,G946);
  nand NAND2_123(G976,G641,G951);
  not NOT_272(G977,G943);
  nand NAND2_124(G980,G924,G962);
  nand NAND2_125(G981,G926,G963);
  nand NAND2_126(G984,G928,G964);
  nand NAND2_127(G987,G930,G967);
  nand NAND2_128(G988,G932,G968);
  nand NAND2_129(G989,G934,G969);
  nand NAND2_130(G993,G936,G970);
  nand NAND2_131(G994,G938,G971);
  not NOT_273(G995,G948);
  nand NAND2_132(G996,G941,G972);
  not NOT_274(G997,G953);
  not NOT_275(G998,G956);
  not NOT_276(G999,G959);
  nand NAND2_133(G1000,G947,G975);
  nand NAND2_134(G1003,G945,G974);
  nand NAND2_135(G1006,G952,G976);
  not NOT_277(G1009,G980);
  not NOT_278(G1012,G988);
  not NOT_279(G1015,G993);
  not NOT_280(G1019,G987);
  nand NAND2_136(G1022,G959,G998);
  nand NAND2_137(G1023,G956,G999);
  not NOT_281(G1024,G977);
  not NOT_282(G1025,G994);
  not NOT_283(G1028,G996);
  not NOT_284(G1031,G989);
  not NOT_285(G1034,G1000);
  not NOT_286(G1035,G1003);
  nand NAND2_138(G1036,G1006,G997);
  not NOT_287(G1037,G1006);
  nand NAND2_139(G1038,G1022,G1023);
  not NOT_288(G1041,G984);
  not NOT_289(G1044,G984);
  not NOT_290(G1047,G989);
  not NOT_291(G1050,G989);
  not NOT_292(G1053,G981);
  not NOT_293(G1056,G981);
  not NOT_294(G1059,G1015);
  not NOT_295(G1062,G1012);
  not NOT_296(G1065,G1025);
  nand NAND2_140(G1066,G953,G1037);
  nand NAND2_141(G1067,G1028,G1024);
  not NOT_297(G1068,G1028);
  not NOT_298(G1069,G1019);
  not NOT_299(G1072,G1019);
  not NOT_300(G1075,G1009);
  not NOT_301(G1078,G1009);
  not NOT_302(G1081,G1012);
  not NOT_303(G1084,G1015);
  not NOT_304(G1087,G1015);
  nand NAND2_142(G1090,G1038,G540);
  not NOT_305(G1091,G1038);
  not NOT_306(G1092,G1041);
  not NOT_307(G1093,G1044);
  nand NAND2_143(G1094,G1047,G784);
  not NOT_308(G1095,G1047);
  nand NAND2_144(G1096,G1050,G786);
  not NOT_309(G1097,G1050);
  not NOT_310(G1098,G1053);
  not NOT_311(G1099,G1056);
  nand NAND2_145(G1100,G1036,G1066);
  nand NAND2_146(G1103,G977,G1068);
  not NOT_312(G1104,G1031);
  not NOT_313(G1107,G1031);
  nand NAND2_147(G1110,G422,G1091);
  not NOT_314(G1111,G1072);
  nand NAND2_148(G1112,G1075,G1092);
  not NOT_315(G1113,G1075);
  nand NAND2_149(G1114,G1078,G1093);
  not NOT_316(G1115,G1078);
  nand NAND2_150(G1116,G675,G1095);
  nand NAND2_151(G1117,G678,G1097);
  not NOT_317(G1118,G1059);
  not NOT_318(G1121,G1059);
  nand NAND2_152(G1124,G1081,G1035);
  not NOT_319(G1125,G1081);
  nand NAND2_153(G1126,G1067,G1103);
  not NOT_320(G1129,G1084);
  not NOT_321(G1130,G1069);
  not NOT_322(G1131,G1087);
  not NOT_323(G1132,G1062);
  not NOT_324(G1135,G1062);
  nand NAND2_154(G1138,G1100,G995);
  not NOT_325(G1139,G1100);
  nand NAND2_155(G1140,G1090,G1110);
  nand NAND2_156(G1143,G1041,G1113);
  nand NAND2_157(G1144,G1044,G1115);
  nand NAND2_158(G1145,G1094,G1116);
  nand NAND2_159(G1148,G1096,G1117);
  nand NAND2_160(G1151,G1003,G1125);
  not NOT_326(G1152,G1104);
  nand NAND2_161(G1153,G1104,G1129);
  not NOT_327(G1154,G1107);
  nand NAND2_162(G1155,G1107,G1131);
  not NOT_328(G1156,G1121);
  nand NAND2_163(G1157,G948,G1139);
  nand NAND2_164(G1158,G1126,G910);
  not NOT_329(G1159,G1126);
  nand NAND2_165(G1160,G1112,G1143);
  nand NAND2_166(G1163,G1114,G1144);
  not NOT_330(G1166,G1132);
  nand NAND2_167(G1167,G1132,G1098);
  not NOT_331(G1168,G1118);
  not NOT_332(G1169,G1135);
  nand NAND2_168(G1170,G1135,G1099);
  nand NAND2_169(G1171,G1124,G1151);
  nand NAND2_170(G1174,G1084,G1152);
  nand NAND2_171(G1175,G1087,G1154);
  nand NAND2_172(G1176,G1148,G722);
  not NOT_333(G1177,G1148);
  nand NAND2_173(G1178,G1138,G1157);
  nand NAND2_174(G1181,G851,G1159);
  nand NAND2_175(G1182,G1140,G212);
  not NOT_334(G1185,G1145);
  nand NAND2_176(G1186,G1145,G785);
  nand NAND2_177(G1187,G1053,G1166);
  nand NAND2_178(G1188,G1056,G1169);
  nand NAND2_179(G1189,G1174,G1153);
  nand NAND2_180(G1192,G1175,G1155);
  not NOT_335(G1195,G1140);
  nand NAND2_181(G1198,G1163,G965);
  not NOT_336(G1199,G1163);
  nand NAND2_182(G1200,G1160,G966);
  not NOT_337(G1201,G1160);
  nand NAND2_183(G1202,G609,G1177);
  nand NAND2_184(G1203,G1171,G908);
  not NOT_338(G1204,G1171);
  nand NAND2_185(G1205,G1158,G1181);
  nand NAND2_186(G1208,G606,G1185);
  nand NAND2_187(G1209,G1187,G1167);
  nand NAND2_188(G1212,G1188,G1170);
  nand NAND2_189(G1215,G914,G1199);
  nand NAND2_190(G1216,G911,G1201);
  nand NAND2_191(G1217,G1176,G1202);
  nand NAND2_192(G1218,G845,G1204);
  nand NAND2_193(G1219,G1192,G1111);
  not NOT_339(G1220,G1192);
  not NOT_340(G1221,G1195);
  nand NAND2_194(G1222,G1178,G212);
  not NOT_341(G1225,G1189);
  nand NAND2_195(G1226,G1189,G1130);
  not NOT_342(G1227,G1178);
  not NOT_343(G1230,G1182);
  not NOT_344(G1233,G1182);
  nand NAND2_196(G1236,G1186,G1208);
  nand NAND2_197(G1239,G1198,G1215);
  nand NAND2_198(G1240,G1200,G1216);
  nand NAND2_199(G1243,G1212,G1156);
  not NOT_345(G1244,G1212);
  nand NAND2_200(G1245,G1203,G1218);
  nand NAND2_201(G1246,G1072,G1220);
  nand NAND2_202(G1247,G1205,G212);
  not NOT_346(G1250,G1209);
  nand NAND2_203(G1251,G1209,G1168);
  nand NAND2_204(G1252,G1069,G1225);
  not NOT_347(G1253,G1217);
  not NOT_348(G1256,G1205);
  not NOT_349(G1259,G1239);
  nand NAND2_205(G1260,G1121,G1244);
  not NOT_350(G1261,G1245);
  nand NAND2_206(G1262,G1219,G1246);
  not NOT_351(G1263,G1227);
  nand NAND2_207(G1264,G1233,G566);
  not NOT_352(G1265,G1233);
  nand NAND2_208(G1266,G1230,G567);
  not NOT_353(G1267,G1230);
  not NOT_354(G1268,G1236);
  nand NAND2_209(G1269,G1118,G1250);
  not NOT_355(G1270,G1222);
  not NOT_356(G1273,G1222);
  nand NAND2_210(G1276,G1226,G1252);
  nand NAND2_211(G1279,G1243,G1260);
  not NOT_357(G1280,G1253);
  not NOT_358(G1281,G1256);
  nand NAND2_212(G1282,G458,G1265);
  nand NAND2_213(G1283,G455,G1267);
  not NOT_359(G1284,G1240);
  not NOT_360(G1287,G1262);
  not NOT_361(G1290,G1247);
  not NOT_362(G1293,G1247);
  not NOT_363(G1296,G1240);
  nand NAND2_214(G1299,G1251,G1269);
  and AND2_6(G1302,G1259,G380);
  and AND2_7(G1305,G381,G1261);
  nand NAND2_215(G1308,G1273,G564);
  not NOT_364(G1309,G1273);
  nand NAND2_216(G1310,G1270,G565);
  not NOT_365(G1311,G1270);
  nand NAND2_217(G1312,G1264,G1282);
  nand NAND2_218(G1313,G1266,G1283);
  not NOT_366(G1316,G1276);
  not NOT_367(G1317,G1279);
  not NOT_368(G1320,G1284);
  nand NAND2_219(G1321,G1284,G1280);
  not NOT_369(G1322,G1287);
  nand NAND2_220(G1323,G1287,G973);
  nand NAND2_221(G1324,G1293,G859);
  not NOT_370(G1325,G1293);
  nand NAND2_222(G1326,G1290,G860);
  not NOT_371(G1327,G1290);
  nand NAND2_223(G1328,G452,G1309);
  nand NAND2_224(G1329,G449,G1311);
  not NOT_372(G1330,G1312);
  not NOT_373(G1331,G1296);
  nand NAND2_225(G1332,G1296,G1268);
  not NOT_374(G1333,G1299);
  nand NAND2_226(G1334,G1299,G1065);
  not NOT_375(G1335,G1302);
  not NOT_376(G1336,G1305);
  nand NAND2_227(G1337,G1253,G1320);
  not NOT_377(G1338,G1317);
  nand NAND2_228(G1339,G1317,G1034);
  nand NAND2_229(G1340,G921,G1322);
  nand NAND2_230(G1341,G828,G1325);
  nand NAND2_231(G1342,G825,G1327);
  nand NAND2_232(G1343,G1308,G1328);
  nand NAND2_233(G1344,G1310,G1329);
  not NOT_378(G1347,G1313);
  not NOT_379(G1350,G1313);
  nand NAND2_234(G1353,G1236,G1331);
  nand NAND2_235(G1354,G1025,G1333);
  nand NAND2_236(G1355,G1337,G1321);
  nand NAND2_237(G1356,G1000,G1338);
  nand NAND2_238(G1357,G1340,G1323);
  nand NAND2_239(G1358,G1324,G1341);
  nand NAND2_240(G1359,G1326,G1342);
  not NOT_380(G1362,G1343);
  nand NAND2_241(G1363,G1353,G1332);
  nand NAND2_242(G1366,G1354,G1334);
  not NOT_381(G1369,G1355);
  nand NAND2_243(G1370,G1356,G1339);
  nand NAND2_244(G1371,G1357,G212);
  not NOT_382(G1374,G1358);
  not NOT_383(G1375,G1344);
  not NOT_384(G1378,G1344);
  not NOT_385(G1381,G1363);
  not NOT_386(G1382,G1366);
  nand NAND2_245(G1383,G1369,G212);
  nand NAND2_246(G1386,G1370,G212);
  not NOT_387(G1389,G1359);
  not NOT_388(G1392,G1359);
  and AND2_8(G1395,G1347,G1375);
  and AND2_9(G1410,G1350,G1375);
  and AND2_10(G1420,G1347,G1378);
  and AND2_11(G1434,G1350,G1378);
  not NOT_389(G1439,G1371);
  not NOT_390(G1442,G1371);
  not NOT_391(G1445,G1383);
  not NOT_392(G1448,G1383);
  not NOT_393(G1451,G1386);
  not NOT_394(G1454,G1386);
  nand NAND2_247(G1457,G1442,G562);
  not NOT_395(G1458,G1442);
  nand NAND2_248(G1459,G1439,G563);
  not NOT_396(G1460,G1439);
  nand NAND2_249(G1461,G1448,G857);
  not NOT_397(G1462,G1448);
  nand NAND2_250(G1463,G1445,G858);
  not NOT_398(G1464,G1445);
  nand NAND2_251(G1465,G1454,G560);
  not NOT_399(G1466,G1454);
  nand NAND2_252(G1467,G1451,G561);
  not NOT_400(G1468,G1451);
  nand NAND2_253(G1469,G446,G1458);
  nand NAND2_254(G1470,G443,G1460);
  nand NAND2_255(G1471,G822,G1462);
  nand NAND2_256(G1472,G819,G1464);
  nand NAND2_257(G1473,G440,G1466);
  nand NAND2_258(G1474,G437,G1468);
  nand NAND2_259(G1475,G1457,G1469);
  nand NAND2_260(G1476,G1459,G1470);
  nand NAND2_261(G1479,G1461,G1471);
  nand NAND2_262(G1480,G1463,G1472);
  nand NAND2_263(G1483,G1465,G1473);
  nand NAND2_264(G1484,G1467,G1474);
  not NOT_401(G1487,G1475);
  not NOT_402(G1488,G1479);
  not NOT_403(G1489,G1483);
  not NOT_404(G1490,G1476);
  not NOT_405(G1493,G1476);
  not NOT_406(G1496,G1480);
  and AND2_12(G1499,G731,G1480);
  not NOT_407(G1502,G1484);
  and AND2_13(G1505,G735,G1484);
  nand NAND8_0(G1508,G1374,G1330,G1362,G1487,G546,G1489,G1488,G550);
  not NOT_408(G1511,G1499);
  not NOT_409(G1522,G1499);
  not NOT_410(G1538,G1505);
  not NOT_411(G1549,G1505);
  and AND2_14(G1563,G1389,G1490);
  and AND2_15(G1576,G1392,G1490);
  and AND2_16(G1584,G1389,G1493);
  and AND2_17(G1598,G1392,G1493);
  and AND4_0(G1607,G260,G1508,G235,G235);
  and AND2_18(G1608,G730,G1496);
  and AND2_19(G1609,G731,G1496);
  and AND2_20(G1624,G734,G1502);
  and AND2_21(G1625,G735,G1502);
  nand NAND5_0(G1642,G1511,G1538,G1584,G1395,G738);
  nand NAND5_1(G1645,G1511,G1538,G1563,G1420,G738);
  nand NAND5_2(G1648,G1511,G1538,G1563,G1410,G738);
  nand NAND5_3(G1651,G1511,G1538,G1576,G1395,G738);
  nand NAND5_4(G1654,G1522,G1538,G1598,G1410,G755);
  nand NAND5_5(G1657,G1522,G1549,G1584,G1434,G755);
  nand NAND5_6(G1660,G1522,G1549,G1598,G1420,G755);
  and AND5_0(G1663,G1511,G1538,G1584,G1395,G738);
  and AND5_1(G1666,G1511,G1538,G1563,G1420,G738);
  and AND5_2(G1669,G1511,G1538,G1563,G1410,G738);
  and AND5_3(G1672,G1511,G1538,G1576,G1395,G738);
  and AND5_4(G1675,G1522,G1538,G1598,G1410,G755);
  and AND5_5(G1678,G1522,G1549,G1584,G1434,G755);
  and AND5_6(G1681,G1522,G1549,G1598,G1420,G755);
  nand NAND5_7(G1684,G1511,G1625,G1584,G1420,G738);
  nand NAND5_8(G1687,G1522,G1625,G1584,G1410,G738);
  nand NAND5_9(G1690,G1522,G1625,G1598,G1395,G738);
  nand NAND5_10(G1693,G1522,G1625,G1563,G1434,G738);
  nand NAND5_11(G1696,G1522,G1625,G1576,G1420,G755);
  nand NAND5_12(G1699,G1609,G1549,G1584,G1420,G755);
  nand NAND5_13(G1702,G1609,G1549,G1584,G1410,G755);
  nand NAND5_14(G1705,G1609,G1549,G1598,G1395,G755);
  nand NAND5_15(G1708,G1609,G1549,G1576,G1420,G755);
  nand NAND5_16(G1711,G1522,G1625,G1563,G1395,G573);
  nand NAND5_17(G1712,G1609,G1549,G1563,G1395,G573);
  nand NAND5_18(G1713,G1609,G1625,G1584,G1395,G573);
  nand NAND5_19(G1714,G1609,G1625,G1563,G1420,G573);
  nand NAND5_20(G1715,G1609,G1625,G1563,G1410,G573);
  nand NAND5_21(G1716,G1609,G1625,G1576,G1395,G573);
  nand NAND5_22(G1717,G1609,G1624,G1563,G1395,G573);
  nand NAND5_23(G1718,G1608,G1625,G1563,G1395,G573);
  and AND5_7(G1719,G1511,G1625,G1584,G1420,G738);
  and AND5_8(G1722,G1522,G1625,G1584,G1410,G738);
  and AND5_9(G1725,G1522,G1625,G1598,G1395,G738);
  and AND5_10(G1728,G1522,G1625,G1563,G1434,G738);
  and AND5_11(G1731,G1522,G1625,G1576,G1420,G755);
  and AND5_12(G1734,G1609,G1549,G1584,G1420,G755);
  and AND5_13(G1737,G1609,G1549,G1584,G1410,G755);
  and AND5_14(G1740,G1609,G1549,G1598,G1395,G755);
  and AND5_15(G1743,G1609,G1549,G1576,G1420,G755);
  nand NAND2_265(G1746,G1663,G313);
  not NOT_412(G1747,G1663);
  nand NAND2_266(G1748,G1666,G314);
  not NOT_413(G1749,G1666);
  nand NAND2_267(G1750,G1669,G315);
  not NOT_414(G1751,G1669);
  nand NAND2_268(G1752,G1672,G316);
  not NOT_415(G1753,G1672);
  nand NAND2_269(G1754,G1675,G322);
  not NOT_416(G1755,G1675);
  nand NAND2_270(G1756,G1678,G327);
  not NOT_417(G1757,G1678);
  nand NAND2_271(G1758,G1681,G328);
  not NOT_418(G1759,G1681);
  and AND8_0(G1760,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718);
  nand NAND2_272(G1761,G265,G1747);
  nand NAND2_273(G1762,G268,G1749);
  nand NAND2_274(G1763,G271,G1751);
  nand NAND2_275(G1764,G274,G1753);
  nand NAND2_276(G1765,G1719,G317);
  not NOT_419(G1766,G1719);
  nand NAND2_277(G1767,G1722,G318);
  not NOT_420(G1768,G1722);
  nand NAND2_278(G1769,G1725,G319);
  not NOT_421(G1770,G1725);
  nand NAND2_279(G1771,G1728,G320);
  not NOT_422(G1772,G1728);
  nand NAND2_280(G1773,G1731,G321);
  not NOT_423(G1774,G1731);
  nand NAND2_281(G1775,G292,G1755);
  nand NAND2_282(G1776,G1734,G323);
  not NOT_424(G1777,G1734);
  nand NAND2_283(G1778,G1737,G324);
  not NOT_425(G1779,G1737);
  nand NAND2_284(G1780,G1740,G325);
  not NOT_426(G1781,G1740);
  nand NAND2_285(G1782,G1743,G326);
  not NOT_427(G1783,G1743);
  nand NAND2_286(G1784,G307,G1757);
  nand NAND2_287(G1785,G310,G1759);
  nand NAND8_1(G1786,G1642,G1645,G1648,G1651,G1684,G1687,G1690,G1693);
  nand NAND8_2(G1787,G1696,G1654,G1699,G1702,G1705,G1708,G1657,G1660);
  and AND8_1(G1788,G1642,G1645,G1648,G1651,G1684,G1687,G1690,G1693);
  and AND8_2(G1791,G1696,G1654,G1699,G1702,G1705,G1708,G1657,G1660);
  nand NAND2_288(G1794,G277,G1766);
  nand NAND2_289(G1795,G280,G1768);
  nand NAND2_290(G1796,G283,G1770);
  nand NAND2_291(G1797,G286,G1772);
  nand NAND2_292(G1798,G289,G1774);
  nand NAND2_293(G1799,G295,G1777);
  nand NAND2_294(G1800,G298,G1779);
  nand NAND2_295(G1801,G301,G1781);
  nand NAND2_296(G1802,G304,G1783);
  and AND2_22(G1803,G1786,G197);
  and AND2_23(G1806,G1787,G198);
  and AND3_5(G1809,G1788,G1791,G1760);
  nand NAND2_297(G1810,G1788,G1791);
  and AND4_1(G1817,G260,G1508,G32,G1809);
  nand NAND2_298(G1818,G1803,G1335);
  not NOT_428(G1819,G1803);
  nand NAND2_299(G1820,G1806,G1336);
  not NOT_429(G1821,G1806);
  and AND3_6(G1822,G544,G205,G1810);
  and AND3_7(G1825,G25,G205,G1810);
  and AND3_8(G1828,G27,G205,G1810);
  and AND3_9(G1831,G28,G205,G1810);
  and AND3_10(G1834,G545,G205,G1810);
  nand NAND2_300(G1837,G1302,G1819);
  nand NAND2_301(G1838,G1305,G1821);
  and AND3_11(G1839,G26,G205,G1810);
  nand NAND2_302(G1842,G1818,G1837);
  nand NAND2_303(G1845,G1820,G1838);
  nand NAND2_304(G1848,G1822,G1381);
  nand NAND2_305(G1849,G1825,G1382);
  nand NAND2_306(G1850,G1828,G1263);
  nand NAND2_307(G1851,G1831,G1221);
  nand NAND2_308(G1852,G1834,G1281);
  not NOT_430(G1853,G1822);
  not NOT_431(G1854,G1825);
  not NOT_432(G1855,G1828);
  not NOT_433(G1856,G1831);
  not NOT_434(G1857,G1834);
  not NOT_435(G1858,G1839);
  nand NAND2_309(G1859,G1839,G1316);
  nand NAND2_310(G1860,G1363,G1853);
  nand NAND2_311(G1861,G1366,G1854);
  nand NAND2_312(G1862,G1227,G1855);
  nand NAND2_313(G1863,G1195,G1856);
  nand NAND2_314(G1864,G1256,G1857);
  nand NAND2_315(G1865,G1842,G533);
  not NOT_436(G1866,G1842);
  nand NAND2_316(G1867,G1845,G534);
  not NOT_437(G1868,G1845);
  nand NAND2_317(G1869,G1276,G1858);
  nand NAND2_318(G1870,G1860,G1848);
  nand NAND2_319(G1871,G1861,G1849);
  nand NAND2_320(G1872,G1862,G1850);
  nand NAND2_321(G1873,G1863,G1851);
  nand NAND2_322(G1874,G1864,G1852);
  nand NAND2_323(G1875,G461,G1866);
  nand NAND2_324(G1876,G464,G1868);
  nand NAND2_325(G1877,G1869,G1859);
  nand NAND2_326(G1880,G1877,G940);
  not NOT_438(G1881,G1877);
  nand NAND2_327(G1882,G891,G1881);
  nand NAND2_328(G1883,G1880,G1882);
  nand NAND2_329(G1884,G1746,G1761);
  nand NAND2_330(G1885,G1748,G1762);
  nand NAND2_331(G1886,G1750,G1763);
  nand NAND2_332(G1887,G1752,G1764);
  nand NAND2_333(G1888,G1754,G1775);
  nand NAND2_334(G1889,G1756,G1784);
  nand NAND2_335(G1890,G1758,G1785);
  nand NAND2_336(G1891,G1765,G1794);
  nand NAND2_337(G1892,G1767,G1795);
  nand NAND2_338(G1893,G1769,G1796);
  nand NAND2_339(G1894,G1771,G1797);
  nand NAND2_340(G1895,G1773,G1798);
  nand NAND2_341(G1896,G1776,G1799);
  nand NAND2_342(G1897,G1778,G1800);
  nand NAND2_343(G1898,G1780,G1801);
  nand NAND2_344(G1899,G1782,G1802);
  nor NOR2_0(G1900,G1607,G1817);
  and AND2_24(G1901,G1870,G329);
  and AND2_25(G1902,G330,G1871);
  and AND2_26(G1903,G332,G1872);
  and AND2_27(G1904,G1873,G333);
  and AND2_28(G1905,G334,G1874);
  nand NAND2_345(G1906,G1865,G1875);
  nand NAND2_346(G1907,G1867,G1876);
  and AND2_29(G1908,G1883,G331);

endmodule
