
//Verilog file of module c3540


`timescale 1 ns / 1ns

module c3540_net(G1,
G10,
G11,
G12,
G13,
G14,
G15,
G16,
G17,
G18,
G19,
G2,
G20,
G21,
G22,
G23,
G24,
G25,
G26,
G27,
G28,
G29,
G3,
G30,
G31,
G32,
G33,
G34,
G35,
G3519,
G3520,
G3521,
G3522,
G3523,
G3524,
G3525,
G3526,
G3527,
G3528,
G3529,
G3530,
G3531,
G3532,
G3533,
G3534,
G3535,
G3536,
G3537,
G3538,
G3539,
G3540,
G36,
G37,
G38,
G39,
G4,
G40,
G41,
G42,
G43,
G44,
G45,
G46,
G47,
G48,
G49,
G5,
G50,
G6,
G7,
G8,
G9);
input G1;
input G2;
input G3;
input G4;
input G5;
input G6;
input G7;
input G8;
input G9;
input G10;
input G11;
input G12;
input G13;
input G14;
input G15;
input G16;
input G17;
input G18;
input G19;
input G20;
input G21;
input G22;
input G23;
input G24;
input G25;
input G26;
input G27;
input G28;
input G29;
input G30;
input G31;
input G32;
input G33;
input G34;
input G35;
input G36;
input G37;
input G38;
input G39;
input G40;
input G41;
input G42;
input G43;
input G44;
input G45;
input G46;
input G47;
input G48;
input G49;
input G50;

output G3519;
output G3520;
output G3521;
output G3522;
output G3523;
output G3524;
output G3525;
output G3526;
output G3527;
output G3528;
output G3529;
output G3530;
output G3531;
output G3532;
output G3533;
output G3534;
output G3535;
output G3536;
output G3537;
output G3538;
output G3539;
output G3540;

wire
c3540_wire_1,
c3540_wire_2,
c3540_wire_3,
c3540_wire_4,
c3540_wire_5,
c3540_wire_6,
c3540_wire_7,
c3540_wire_8,
c3540_wire_9,
c3540_wire_10,
c3540_wire_11,
c3540_wire_12,
c3540_wire_13,
c3540_wire_14,
c3540_wire_15,
c3540_wire_16,
c3540_wire_17,
c3540_wire_18,
c3540_wire_19,
c3540_wire_20,
c3540_wire_21,
c3540_wire_22,
c3540_wire_23,
c3540_wire_24,
c3540_wire_25,
c3540_wire_26,
c3540_wire_27,
c3540_wire_28,
c3540_wire_29,
c3540_wire_30,
c3540_wire_31,
c3540_wire_32,
c3540_wire_33,
c3540_wire_34,
c3540_wire_35,
c3540_wire_36,
c3540_wire_37,
c3540_wire_38,
c3540_wire_39,
c3540_wire_40,
c3540_wire_41,
c3540_wire_42,
c3540_wire_43,
c3540_wire_44,
c3540_wire_45,
c3540_wire_46,
c3540_wire_47,
c3540_wire_48,
c3540_wire_49,
c3540_wire_50,
c3540_wire_51,
c3540_wire_52,
c3540_wire_53,
c3540_wire_54,
c3540_wire_55,
c3540_wire_56,
c3540_wire_57,
c3540_wire_58,
c3540_wire_59,
c3540_wire_60,
c3540_wire_61,
c3540_wire_62,
c3540_wire_63,
c3540_wire_64,
c3540_wire_65,
c3540_wire_66,
c3540_wire_67,
c3540_wire_68,
c3540_wire_69,
c3540_wire_70,
c3540_wire_71,
c3540_wire_72,
c3540_wire_73,
c3540_wire_74,
c3540_wire_75,
c3540_wire_76,
c3540_wire_77,
c3540_wire_78,
c3540_wire_79,
c3540_wire_80,
c3540_wire_81,
c3540_wire_82,
c3540_wire_83,
c3540_wire_84,
c3540_wire_85,
c3540_wire_86,
c3540_wire_87,
c3540_wire_88,
c3540_wire_89,
c3540_wire_90,
c3540_wire_91,
c3540_wire_92,
c3540_wire_93,
c3540_wire_94,
c3540_wire_95,
c3540_wire_96,
c3540_wire_97,
c3540_wire_98,
c3540_wire_99,
c3540_wire_100,
c3540_wire_101,
c3540_wire_102,
c3540_wire_103,
c3540_wire_104,
c3540_wire_105,
c3540_wire_106,
c3540_wire_107,
c3540_wire_108,
c3540_wire_109,
c3540_wire_110,
c3540_wire_111,
c3540_wire_112,
c3540_wire_113,
c3540_wire_114,
c3540_wire_115,
c3540_wire_116,
c3540_wire_117,
c3540_wire_118,
c3540_wire_119,
c3540_wire_120,
c3540_wire_121,
c3540_wire_122,
c3540_wire_123,
c3540_wire_124,
c3540_wire_125,
c3540_wire_126,
c3540_wire_127,
c3540_wire_128,
c3540_wire_129,
c3540_wire_130,
c3540_wire_131,
c3540_wire_132,
c3540_wire_133,
c3540_wire_134,
c3540_wire_135,
c3540_wire_136,
c3540_wire_137,
c3540_wire_138,
c3540_wire_139,
c3540_wire_140,
c3540_wire_141,
c3540_wire_142,
c3540_wire_143,
c3540_wire_144,
c3540_wire_145,
c3540_wire_146,
c3540_wire_147,
c3540_wire_148,
c3540_wire_149,
c3540_wire_150,
c3540_wire_151,
c3540_wire_152,
c3540_wire_153,
c3540_wire_154,
c3540_wire_155,
c3540_wire_156,
c3540_wire_157,
c3540_wire_158,
c3540_wire_159,
c3540_wire_160,
c3540_wire_161,
c3540_wire_162,
c3540_wire_163,
c3540_wire_164,
c3540_wire_165,
c3540_wire_166,
c3540_wire_167,
c3540_wire_168,
c3540_wire_169,
c3540_wire_170,
c3540_wire_171,
c3540_wire_172,
c3540_wire_173,
c3540_wire_174,
c3540_wire_175,
c3540_wire_176,
c3540_wire_177,
c3540_wire_178,
c3540_wire_179,
c3540_wire_180,
c3540_wire_181,
c3540_wire_182,
c3540_wire_183,
c3540_wire_184,
c3540_wire_185,
c3540_wire_186,
c3540_wire_187,
c3540_wire_188,
c3540_wire_189,
c3540_wire_190,
c3540_wire_191,
c3540_wire_192,
c3540_wire_193,
c3540_wire_194,
c3540_wire_195,
c3540_wire_196,
c3540_wire_197,
c3540_wire_198,
c3540_wire_199,
c3540_wire_200,
c3540_wire_201,
c3540_wire_202,
c3540_wire_203,
c3540_wire_204,
c3540_wire_205,
c3540_wire_206,
c3540_wire_207,
c3540_wire_208,
c3540_wire_209,
c3540_wire_210,
c3540_wire_211,
c3540_wire_212,
c3540_wire_213,
c3540_wire_214,
c3540_wire_215,
c3540_wire_216,
c3540_wire_217,
c3540_wire_218,
c3540_wire_219,
c3540_wire_220,
c3540_wire_221,
c3540_wire_222,
c3540_wire_223,
c3540_wire_224,
c3540_wire_225,
c3540_wire_226,
c3540_wire_227,
c3540_wire_228,
c3540_wire_229,
c3540_wire_230,
c3540_wire_231,
c3540_wire_232,
c3540_wire_233,
c3540_wire_234,
c3540_wire_235,
c3540_wire_236,
c3540_wire_237,
c3540_wire_238,
c3540_wire_239,
c3540_wire_240,
c3540_wire_241,
c3540_wire_242,
c3540_wire_243,
c3540_wire_244,
c3540_wire_245,
c3540_wire_246,
c3540_wire_247,
c3540_wire_248,
c3540_wire_249,
c3540_wire_250,
c3540_wire_251,
c3540_wire_252,
c3540_wire_253,
c3540_wire_254,
c3540_wire_255,
c3540_wire_256,
c3540_wire_257,
c3540_wire_258,
c3540_wire_259,
c3540_wire_260,
c3540_wire_261,
c3540_wire_262,
c3540_wire_263,
c3540_wire_264,
c3540_wire_265,
c3540_wire_266,
c3540_wire_267,
c3540_wire_268,
c3540_wire_269,
c3540_wire_270,
c3540_wire_271,
c3540_wire_272,
c3540_wire_273,
c3540_wire_274,
c3540_wire_275,
c3540_wire_276,
c3540_wire_277,
c3540_wire_278,
c3540_wire_279,
c3540_wire_280,
c3540_wire_281,
c3540_wire_282,
c3540_wire_283,
c3540_wire_284,
c3540_wire_285,
c3540_wire_286,
c3540_wire_287,
c3540_wire_288,
c3540_wire_289,
c3540_wire_290,
c3540_wire_291,
c3540_wire_292,
c3540_wire_293,
c3540_wire_294,
c3540_wire_295,
c3540_wire_296,
c3540_wire_297,
c3540_wire_298,
c3540_wire_299,
c3540_wire_300,
c3540_wire_301,
c3540_wire_302,
c3540_wire_303,
c3540_wire_304,
c3540_wire_305,
c3540_wire_306,
c3540_wire_307,
c3540_wire_308,
c3540_wire_309,
c3540_wire_310,
c3540_wire_311,
c3540_wire_312,
c3540_wire_313,
c3540_wire_314,
c3540_wire_315,
c3540_wire_316,
c3540_wire_317,
c3540_wire_318,
c3540_wire_319,
c3540_wire_320,
c3540_wire_321,
c3540_wire_322,
c3540_wire_323,
c3540_wire_324,
c3540_wire_325,
c3540_wire_326,
c3540_wire_327,
c3540_wire_328,
c3540_wire_329,
c3540_wire_330,
c3540_wire_331,
c3540_wire_332,
c3540_wire_333,
c3540_wire_334,
c3540_wire_335,
c3540_wire_336,
c3540_wire_337,
c3540_wire_338,
c3540_wire_339,
c3540_wire_340,
c3540_wire_341,
c3540_wire_342,
c3540_wire_343,
c3540_wire_344,
c3540_wire_345,
c3540_wire_346,
c3540_wire_347,
c3540_wire_348,
c3540_wire_349,
c3540_wire_350,
c3540_wire_351,
c3540_wire_352,
c3540_wire_353,
c3540_wire_354,
c3540_wire_355,
c3540_wire_356,
c3540_wire_357,
c3540_wire_358,
c3540_wire_359,
c3540_wire_360,
c3540_wire_361,
c3540_wire_362,
c3540_wire_363,
c3540_wire_364,
c3540_wire_365,
c3540_wire_366,
c3540_wire_367,
c3540_wire_368,
c3540_wire_369,
c3540_wire_370,
c3540_wire_371,
c3540_wire_372,
c3540_wire_373,
c3540_wire_374,
c3540_wire_375,
c3540_wire_376,
c3540_wire_377,
c3540_wire_378,
c3540_wire_379,
c3540_wire_380,
c3540_wire_381,
c3540_wire_382,
c3540_wire_383,
c3540_wire_384,
c3540_wire_385,
c3540_wire_386,
c3540_wire_387,
c3540_wire_388,
c3540_wire_389,
c3540_wire_390,
c3540_wire_391,
c3540_wire_392,
c3540_wire_393,
c3540_wire_394,
c3540_wire_395,
c3540_wire_396,
c3540_wire_397,
c3540_wire_398,
c3540_wire_399,
c3540_wire_400,
c3540_wire_401,
c3540_wire_402,
c3540_wire_403,
c3540_wire_404,
c3540_wire_405,
c3540_wire_406,
c3540_wire_407,
c3540_wire_408,
c3540_wire_409,
c3540_wire_410,
c3540_wire_411,
c3540_wire_412,
c3540_wire_413,
c3540_wire_414,
c3540_wire_415,
c3540_wire_416,
c3540_wire_417,
c3540_wire_418,
c3540_wire_419,
c3540_wire_420,
c3540_wire_421,
c3540_wire_422,
c3540_wire_423,
c3540_wire_424,
c3540_wire_425,
c3540_wire_426,
c3540_wire_427,
c3540_wire_428,
c3540_wire_429,
c3540_wire_430,
c3540_wire_431,
c3540_wire_432,
c3540_wire_433,
c3540_wire_434,
c3540_wire_435,
c3540_wire_436,
c3540_wire_437,
c3540_wire_438,
c3540_wire_439,
c3540_wire_440,
c3540_wire_441,
c3540_wire_442,
c3540_wire_443,
c3540_wire_444,
c3540_wire_445,
c3540_wire_446,
c3540_wire_447,
c3540_wire_448,
c3540_wire_449,
c3540_wire_450,
c3540_wire_451,
c3540_wire_452,
c3540_wire_453,
c3540_wire_454,
c3540_wire_455,
c3540_wire_456,
c3540_wire_457,
c3540_wire_458,
c3540_wire_459,
c3540_wire_460,
c3540_wire_461,
c3540_wire_462,
c3540_wire_463,
c3540_wire_464,
c3540_wire_465,
c3540_wire_466,
c3540_wire_467,
c3540_wire_468,
c3540_wire_469,
c3540_wire_470,
c3540_wire_471,
c3540_wire_472,
c3540_wire_473,
c3540_wire_474,
c3540_wire_475,
c3540_wire_476,
c3540_wire_477,
c3540_wire_478,
c3540_wire_479,
c3540_wire_480,
c3540_wire_481,
c3540_wire_482,
c3540_wire_483,
c3540_wire_484,
c3540_wire_485,
c3540_wire_486,
c3540_wire_487,
c3540_wire_488,
c3540_wire_489,
c3540_wire_490,
c3540_wire_491,
c3540_wire_492,
c3540_wire_493,
c3540_wire_494,
c3540_wire_495,
c3540_wire_496,
c3540_wire_497,
c3540_wire_498,
c3540_wire_499,
c3540_wire_500,
c3540_wire_501,
c3540_wire_502,
c3540_wire_503,
c3540_wire_504,
c3540_wire_505,
c3540_wire_506,
c3540_wire_507,
c3540_wire_508,
c3540_wire_509,
c3540_wire_510,
c3540_wire_511,
c3540_wire_512,
c3540_wire_513,
c3540_wire_514,
c3540_wire_515,
c3540_wire_516,
c3540_wire_517,
c3540_wire_518,
c3540_wire_519,
c3540_wire_520,
c3540_wire_521,
c3540_wire_522,
c3540_wire_523,
c3540_wire_524,
c3540_wire_525,
c3540_wire_526,
c3540_wire_527,
c3540_wire_528,
c3540_wire_529,
c3540_wire_530,
c3540_wire_531,
c3540_wire_532,
c3540_wire_533,
c3540_wire_534,
c3540_wire_535,
c3540_wire_536,
c3540_wire_537,
c3540_wire_538,
c3540_wire_539,
c3540_wire_540,
c3540_wire_541,
c3540_wire_542,
c3540_wire_543,
c3540_wire_544,
c3540_wire_545,
c3540_wire_546,
c3540_wire_547,
c3540_wire_548,
c3540_wire_549,
c3540_wire_550,
c3540_wire_551,
c3540_wire_552,
c3540_wire_553,
c3540_wire_554,
c3540_wire_555,
c3540_wire_556,
c3540_wire_557,
c3540_wire_558,
c3540_wire_559,
c3540_wire_560,
c3540_wire_561,
c3540_wire_562,
c3540_wire_563,
c3540_wire_564,
c3540_wire_565,
c3540_wire_566,
c3540_wire_567,
c3540_wire_568,
c3540_wire_569,
c3540_wire_570,
c3540_wire_571,
c3540_wire_572,
c3540_wire_573,
c3540_wire_574,
c3540_wire_575,
c3540_wire_576,
c3540_wire_577,
c3540_wire_578,
c3540_wire_579,
c3540_wire_580,
c3540_wire_581,
c3540_wire_582,
c3540_wire_583,
c3540_wire_584,
c3540_wire_585,
c3540_wire_586,
c3540_wire_587,
c3540_wire_588,
c3540_wire_589,
c3540_wire_590,
c3540_wire_591,
c3540_wire_592,
c3540_wire_593,
c3540_wire_594,
c3540_wire_595,
c3540_wire_596,
c3540_wire_597,
c3540_wire_598,
c3540_wire_599,
c3540_wire_600,
c3540_wire_601,
c3540_wire_602,
c3540_wire_603,
c3540_wire_604,
c3540_wire_605,
c3540_wire_606,
c3540_wire_607,
c3540_wire_608,
c3540_wire_609,
c3540_wire_610,
c3540_wire_611,
c3540_wire_612,
c3540_wire_613,
c3540_wire_614,
c3540_wire_615,
c3540_wire_616,
c3540_wire_617,
c3540_wire_618,
c3540_wire_619,
c3540_wire_620,
c3540_wire_621,
c3540_wire_622,
c3540_wire_623,
c3540_wire_624,
c3540_wire_625,
c3540_wire_626,
c3540_wire_627,
c3540_wire_628,
c3540_wire_629,
c3540_wire_630,
c3540_wire_631,
c3540_wire_632,
c3540_wire_633,
c3540_wire_634,
c3540_wire_635,
c3540_wire_636,
c3540_wire_637,
c3540_wire_638,
c3540_wire_639,
c3540_wire_640,
c3540_wire_641,
c3540_wire_642,
c3540_wire_643,
c3540_wire_644,
c3540_wire_645,
c3540_wire_646,
c3540_wire_647,
c3540_wire_648,
c3540_wire_649,
c3540_wire_650,
c3540_wire_651,
c3540_wire_652,
c3540_wire_653,
c3540_wire_654,
c3540_wire_655,
c3540_wire_656,
c3540_wire_657,
c3540_wire_658,
c3540_wire_659,
c3540_wire_660,
c3540_wire_661,
c3540_wire_662,
c3540_wire_663,
c3540_wire_664,
c3540_wire_665,
c3540_wire_666,
c3540_wire_667,
c3540_wire_668,
c3540_wire_669,
c3540_wire_670,
c3540_wire_671,
c3540_wire_672,
c3540_wire_673,
c3540_wire_674,
c3540_wire_675,
c3540_wire_676,
c3540_wire_677,
c3540_wire_678,
c3540_wire_679,
c3540_wire_680,
c3540_wire_681,
c3540_wire_682,
c3540_wire_683,
c3540_wire_684,
c3540_wire_685,
c3540_wire_686,
c3540_wire_687,
c3540_wire_688,
c3540_wire_689,
c3540_wire_690,
c3540_wire_691,
c3540_wire_692,
c3540_wire_693,
c3540_wire_694,
c3540_wire_695,
c3540_wire_696,
c3540_wire_697,
c3540_wire_698,
c3540_wire_699,
c3540_wire_700,
c3540_wire_701,
c3540_wire_702,
c3540_wire_703,
c3540_wire_704,
c3540_wire_705,
c3540_wire_706,
c3540_wire_707,
c3540_wire_708,
c3540_wire_709,
c3540_wire_710,
c3540_wire_711,
c3540_wire_712,
c3540_wire_713,
c3540_wire_714,
c3540_wire_715,
c3540_wire_716,
c3540_wire_717,
c3540_wire_718,
c3540_wire_719,
c3540_wire_720,
c3540_wire_721,
c3540_wire_722,
c3540_wire_723,
c3540_wire_724,
c3540_wire_725,
c3540_wire_726,
c3540_wire_727,
c3540_wire_728,
c3540_wire_729,
c3540_wire_730,
c3540_wire_731,
c3540_wire_732,
c3540_wire_733,
c3540_wire_734,
c3540_wire_735,
c3540_wire_736,
c3540_wire_737,
c3540_wire_738,
c3540_wire_739,
c3540_wire_740,
c3540_wire_741,
c3540_wire_742,
c3540_wire_743,
c3540_wire_744,
c3540_wire_745,
c3540_wire_746,
c3540_wire_747,
c3540_wire_748,
c3540_wire_749,
c3540_wire_750,
c3540_wire_751,
c3540_wire_752,
c3540_wire_753,
c3540_wire_754,
c3540_wire_755,
c3540_wire_756,
c3540_wire_757,
c3540_wire_758,
c3540_wire_759,
c3540_wire_760,
c3540_wire_761,
c3540_wire_762,
c3540_wire_763,
c3540_wire_764,
c3540_wire_765,
c3540_wire_766,
c3540_wire_767,
c3540_wire_768,
c3540_wire_769,
c3540_wire_770,
c3540_wire_771,
c3540_wire_772,
c3540_wire_773,
c3540_wire_774,
c3540_wire_775,
c3540_wire_776,
c3540_wire_777,
c3540_wire_778,
c3540_wire_779,
c3540_wire_780,
c3540_wire_781,
c3540_wire_782,
c3540_wire_783,
c3540_wire_784,
c3540_wire_785,
c3540_wire_786,
c3540_wire_787,
c3540_wire_788,
c3540_wire_789,
c3540_wire_790,
c3540_wire_791,
c3540_wire_792,
c3540_wire_793,
c3540_wire_794,
c3540_wire_795,
c3540_wire_796,
c3540_wire_797,
c3540_wire_798,
c3540_wire_799,
c3540_wire_800,
c3540_wire_801,
c3540_wire_802,
c3540_wire_803,
c3540_wire_804,
c3540_wire_805,
c3540_wire_806,
c3540_wire_807,
c3540_wire_808,
c3540_wire_809,
c3540_wire_810,
c3540_wire_811,
c3540_wire_812,
c3540_wire_813,
c3540_wire_814,
c3540_wire_815,
c3540_wire_816,
c3540_wire_817,
c3540_wire_818,
c3540_wire_819,
c3540_wire_820,
c3540_wire_821,
c3540_wire_822,
c3540_wire_823,
c3540_wire_824,
c3540_wire_825,
c3540_wire_826,
c3540_wire_827,
c3540_wire_828,
c3540_wire_829,
c3540_wire_830,
c3540_wire_831,
c3540_wire_832,
c3540_wire_833,
c3540_wire_834,
c3540_wire_835,
c3540_wire_836,
c3540_wire_837,
c3540_wire_838,
c3540_wire_839,
c3540_wire_840,
c3540_wire_841,
c3540_wire_842,
c3540_wire_843,
c3540_wire_844,
c3540_wire_845,
c3540_wire_846,
c3540_wire_847,
c3540_wire_848,
c3540_wire_849,
c3540_wire_850,
c3540_wire_851,
c3540_wire_852,
c3540_wire_853,
c3540_wire_854,
c3540_wire_855,
c3540_wire_856,
c3540_wire_857,
c3540_wire_858,
c3540_wire_859,
c3540_wire_860,
c3540_wire_861,
c3540_wire_862,
c3540_wire_863,
c3540_wire_864,
c3540_wire_865,
c3540_wire_866,
c3540_wire_867,
c3540_wire_868,
c3540_wire_869,
c3540_wire_870,
c3540_wire_871,
c3540_wire_872,
c3540_wire_873,
c3540_wire_874,
c3540_wire_875,
c3540_wire_876,
c3540_wire_877,
c3540_wire_878,
c3540_wire_879,
c3540_wire_880,
c3540_wire_881,
c3540_wire_882,
c3540_wire_883,
c3540_wire_884,
c3540_wire_885,
c3540_wire_886,
c3540_wire_887,
c3540_wire_888,
c3540_wire_889,
c3540_wire_890,
c3540_wire_891,
c3540_wire_892,
c3540_wire_893,
c3540_wire_894,
c3540_wire_895,
c3540_wire_896,
c3540_wire_897,
c3540_wire_898,
c3540_wire_899,
c3540_wire_900,
c3540_wire_901,
c3540_wire_902,
c3540_wire_903,
c3540_wire_904,
c3540_wire_905,
c3540_wire_906,
c3540_wire_907,
c3540_wire_908,
c3540_wire_909,
c3540_wire_910,
c3540_wire_911,
c3540_wire_912,
c3540_wire_913,
c3540_wire_914,
c3540_wire_915,
c3540_wire_916,
c3540_wire_917,
c3540_wire_918,
c3540_wire_919,
c3540_wire_920,
c3540_wire_921,
c3540_wire_922,
c3540_wire_923,
c3540_wire_924,
c3540_wire_925,
c3540_wire_926,
c3540_wire_927,
c3540_wire_928,
c3540_wire_929,
c3540_wire_930,
c3540_wire_931,
c3540_wire_932,
c3540_wire_933,
c3540_wire_934,
c3540_wire_935,
c3540_wire_936,
c3540_wire_937,
c3540_wire_938,
c3540_wire_939,
c3540_wire_940,
c3540_wire_941,
c3540_wire_942,
c3540_wire_943,
c3540_wire_944,
c3540_wire_945,
c3540_wire_946,
c3540_wire_947,
c3540_wire_948,
c3540_wire_949,
c3540_wire_950,
c3540_wire_951,
c3540_wire_952,
c3540_wire_953,
c3540_wire_954,
c3540_wire_955,
c3540_wire_956,
c3540_wire_957,
c3540_wire_958,
c3540_wire_959,
c3540_wire_960,
c3540_wire_961,
c3540_wire_962,
c3540_wire_963,
c3540_wire_964,
c3540_wire_965,
c3540_wire_966,
c3540_wire_967,
c3540_wire_968,
c3540_wire_969,
c3540_wire_970,
c3540_wire_971,
c3540_wire_972,
c3540_wire_973,
c3540_wire_974,
c3540_wire_975,
c3540_wire_976,
c3540_wire_977,
c3540_wire_978,
c3540_wire_979,
c3540_wire_980,
c3540_wire_981,
c3540_wire_982,
c3540_wire_983,
c3540_wire_984,
c3540_wire_985,
c3540_wire_986,
c3540_wire_987,
c3540_wire_988,
c3540_wire_989,
c3540_wire_990,
c3540_wire_991,
c3540_wire_992,
c3540_wire_993,
c3540_wire_994,
c3540_wire_995,
c3540_wire_996,
c3540_wire_997,
c3540_wire_998,
c3540_wire_999,
c3540_wire_1000,
c3540_wire_1001,
c3540_wire_1002,
c3540_wire_1003,
c3540_wire_1004,
c3540_wire_1005,
c3540_wire_1006,
c3540_wire_1007,
c3540_wire_1008,
c3540_wire_1009,
c3540_wire_1010,
c3540_wire_1011,
c3540_wire_1012,
c3540_wire_1013,
c3540_wire_1014,
c3540_wire_1015,
c3540_wire_1016,
c3540_wire_1017,
c3540_wire_1018,
c3540_wire_1019,
c3540_wire_1020,
c3540_wire_1021,
c3540_wire_1022,
c3540_wire_1023,
c3540_wire_1024,
c3540_wire_1025,
c3540_wire_1026,
c3540_wire_1027,
c3540_wire_1028,
c3540_wire_1029,
c3540_wire_1030,
c3540_wire_1031,
c3540_wire_1032,
c3540_wire_1033,
c3540_wire_1034,
c3540_wire_1035,
c3540_wire_1036,
c3540_wire_1037,
c3540_wire_1038,
c3540_wire_1039,
c3540_wire_1040,
c3540_wire_1041,
c3540_wire_1042,
c3540_wire_1043,
c3540_wire_1044,
c3540_wire_1045,
c3540_wire_1046,
c3540_wire_1047,
c3540_wire_1048,
c3540_wire_1049,
c3540_wire_1050,
c3540_wire_1051,
c3540_wire_1052,
c3540_wire_1053,
c3540_wire_1054,
c3540_wire_1055,
c3540_wire_1056,
c3540_wire_1057,
c3540_wire_1058,
c3540_wire_1059,
c3540_wire_1060,
c3540_wire_1061,
c3540_wire_1062,
c3540_wire_1063,
c3540_wire_1064,
c3540_wire_1065,
c3540_wire_1066,
c3540_wire_1067,
c3540_wire_1068,
c3540_wire_1069,
c3540_wire_1070,
c3540_wire_1071,
c3540_wire_1072,
c3540_wire_1073,
c3540_wire_1074,
c3540_wire_1075,
c3540_wire_1076,
c3540_wire_1077,
c3540_wire_1078,
c3540_wire_1079,
c3540_wire_1080,
c3540_wire_1081,
c3540_wire_1082,
c3540_wire_1083,
c3540_wire_1084,
c3540_wire_1085,
c3540_wire_1086,
c3540_wire_1087,
c3540_wire_1088,
c3540_wire_1089,
c3540_wire_1090,
c3540_wire_1091,
c3540_wire_1092,
c3540_wire_1093,
c3540_wire_1094,
c3540_wire_1095,
c3540_wire_1096,
c3540_wire_1097,
c3540_wire_1098,
c3540_wire_1099,
c3540_wire_1100,
c3540_wire_1101,
c3540_wire_1102,
c3540_wire_1103,
c3540_wire_1104,
c3540_wire_1105,
c3540_wire_1106,
c3540_wire_1107,
c3540_wire_1108,
c3540_wire_1109,
c3540_wire_1110,
c3540_wire_1111,
c3540_wire_1112,
c3540_wire_1113,
c3540_wire_1114,
c3540_wire_1115,
c3540_wire_1116,
c3540_wire_1117,
c3540_wire_1118,
c3540_wire_1119,
c3540_wire_1120,
c3540_wire_1121,
c3540_wire_1122,
c3540_wire_1123,
c3540_wire_1124,
c3540_wire_1125,
c3540_wire_1126,
c3540_wire_1127,
c3540_wire_1128,
c3540_wire_1129,
c3540_wire_1130,
c3540_wire_1131,
c3540_wire_1132,
c3540_wire_1133,
c3540_wire_1134,
c3540_wire_1135,
c3540_wire_1136,
c3540_wire_1137,
c3540_wire_1138,
c3540_wire_1139,
c3540_wire_1140,
c3540_wire_1141,
c3540_wire_1142,
c3540_wire_1143,
c3540_wire_1144,
c3540_wire_1145,
c3540_wire_1146,
c3540_wire_1147,
c3540_wire_1148,
c3540_wire_1149,
c3540_wire_1150,
c3540_wire_1151,
c3540_wire_1152,
c3540_wire_1153,
c3540_wire_1154,
c3540_wire_1155,
c3540_wire_1156,
c3540_wire_1157,
c3540_wire_1158,
c3540_wire_1159,
c3540_wire_1160,
c3540_wire_1161,
c3540_wire_1162,
c3540_wire_1163,
c3540_wire_1164,
c3540_wire_1165,
c3540_wire_1166,
c3540_wire_1167,
c3540_wire_1168,
c3540_wire_1169,
c3540_wire_1170,
c3540_wire_1171,
c3540_wire_1172,
c3540_wire_1173,
c3540_wire_1174,
c3540_wire_1175,
c3540_wire_1176,
c3540_wire_1177,
c3540_wire_1178,
c3540_wire_1179,
c3540_wire_1180,
c3540_wire_1181,
c3540_wire_1182,
c3540_wire_1183,
c3540_wire_1184,
c3540_wire_1185,
c3540_wire_1186,
c3540_wire_1187,
c3540_wire_1188,
c3540_wire_1189,
c3540_wire_1190,
c3540_wire_1191,
c3540_wire_1192,
c3540_wire_1193,
c3540_wire_1194,
c3540_wire_1195,
c3540_wire_1196,
c3540_wire_1197,
c3540_wire_1198,
c3540_wire_1199,
c3540_wire_1200,
c3540_wire_1201,
c3540_wire_1202,
c3540_wire_1203,
c3540_wire_1204,
c3540_wire_1205,
c3540_wire_1206,
c3540_wire_1207,
c3540_wire_1208,
c3540_wire_1209,
c3540_wire_1210,
c3540_wire_1211,
c3540_wire_1212,
c3540_wire_1213,
c3540_wire_1214,
c3540_wire_1215,
c3540_wire_1216,
c3540_wire_1217,
c3540_wire_1218,
c3540_wire_1219,
c3540_wire_1220,
c3540_wire_1221,
c3540_wire_1222,
c3540_wire_1223,
c3540_wire_1224,
c3540_wire_1225,
c3540_wire_1226,
c3540_wire_1227,
c3540_wire_1_0,
c3540_wire_1_1,
c3540_wire_1_2,
c3540_wire_1_3,
c3540_wire_1_4,
c3540_wire_1_5,
c3540_wire_1_6,
c3540_wire_1_7,
c3540_wire_1_8,
c3540_wire_1_9,
c3540_wire_1_10,
c3540_wire_1_11,
c3540_wire_1_12,
c3540_wire_1_13,
c3540_wire_1_14,
c3540_wire_1_15,
c3540_wire_1_16,
c3540_wire_1_17,
c3540_wire_1_18,
c3540_wire_1_19,
c3540_wire_1_20,
c3540_wire_1_21,
c3540_wire_1_22,
c3540_wire_1_23,
c3540_wire_1_24,
c3540_wire_1_25,
c3540_wire_1_26,
c3540_wire_1_27,
c3540_wire_2_0,
c3540_wire_2_1,
c3540_wire_2_2,
c3540_wire_2_3,
c3540_wire_2_4,
c3540_wire_2_5,
c3540_wire_2_6,
c3540_wire_2_7,
c3540_wire_2_8,
c3540_wire_2_9,
c3540_wire_2_10,
c3540_wire_2_11,
c3540_wire_2_12,
c3540_wire_2_13,
c3540_wire_2_14,
c3540_wire_2_15,
c3540_wire_2_16,
c3540_wire_11_0,
c3540_wire_11_1,
c3540_wire_30_0,
c3540_wire_30_1,
c3540_wire_35_0,
c3540_wire_35_1,
c3540_wire_35_2,
c3540_wire_35_3,
c3540_wire_35_4,
c3540_wire_35_5,
c3540_wire_35_6,
c3540_wire_35_7,
c3540_wire_35_8,
c3540_wire_39_0,
c3540_wire_39_1,
c3540_wire_39_2,
c3540_wire_39_3,
c3540_wire_39_4,
c3540_wire_39_5,
c3540_wire_40_0,
c3540_wire_40_1,
c3540_wire_40_2,
c3540_wire_40_3,
c3540_wire_40_4,
c3540_wire_40_5,
c3540_wire_40_6,
c3540_wire_40_7,
c3540_wire_40_8,
c3540_wire_40_9,
c3540_wire_40_10,
c3540_wire_40_11,
c3540_wire_40_12,
c3540_wire_40_13,
c3540_wire_40_14,
c3540_wire_40_15,
c3540_wire_40_16,
c3540_wire_40_17,
c3540_wire_40_18,
c3540_wire_40_19,
c3540_wire_40_20,
c3540_wire_40_21,
c3540_wire_40_22,
c3540_wire_5_0,
c3540_wire_5_1,
c3540_wire_5_2,
c3540_wire_5_3,
c3540_wire_5_4,
c3540_wire_5_5,
c3540_wire_5_6,
c3540_wire_5_7,
c3540_wire_5_8,
c3540_wire_5_9,
c3540_wire_5_10,
c3540_wire_5_11,
c3540_wire_5_12,
c3540_wire_5_13,
c3540_wire_5_14,
c3540_wire_5_15,
c3540_wire_93_0,
c3540_wire_93_1,
c3540_wire_93_2,
c3540_wire_99_0,
c3540_wire_99_1,
c3540_wire_99_2,
c3540_wire_99_3,
c3540_wire_99_4,
c3540_wire_99_5,
c3540_wire_99_6,
c3540_wire_99_7,
c3540_wire_99_8,
c3540_wire_99_9,
c3540_wire_99_10,
c3540_wire_99_11,
c3540_wire_99_12,
c3540_wire_99_13,
c3540_wire_99_14,
c3540_wire_99_15,
c3540_wire_99_16,
c3540_wire_112_0,
c3540_wire_112_1,
c3540_wire_117_0,
c3540_wire_117_1,
c3540_wire_119_0,
c3540_wire_119_1,
c3540_wire_125_0,
c3540_wire_125_1,
c3540_wire_123_0,
c3540_wire_123_1,
c3540_wire_123_2,
c3540_wire_123_3,
c3540_wire_123_4,
c3540_wire_123_5,
c3540_wire_123_6,
c3540_wire_123_7,
c3540_wire_123_8,
c3540_wire_123_9,
c3540_wire_123_10,
c3540_wire_123_11,
c3540_wire_123_12,
c3540_wire_123_13,
c3540_wire_123_14,
c3540_wire_123_15,
c3540_wire_153_0,
c3540_wire_153_1,
c3540_wire_153_2,
c3540_wire_153_3,
c3540_wire_153_4,
c3540_wire_153_5,
c3540_wire_153_6,
c3540_wire_153_7,
c3540_wire_155_0,
c3540_wire_155_1,
c3540_wire_155_2,
c3540_wire_155_3,
c3540_wire_155_4,
c3540_wire_155_5,
c3540_wire_155_6,
c3540_wire_155_7,
c3540_wire_155_8,
c3540_wire_155_9,
c3540_wire_155_10,
c3540_wire_155_11,
c3540_wire_155_12,
c3540_wire_155_13,
c3540_wire_155_14,
c3540_wire_155_15,
c3540_wire_157_0,
c3540_wire_157_1,
c3540_wire_157_2,
c3540_wire_157_3,
c3540_wire_157_4,
c3540_wire_157_5,
c3540_wire_157_6,
c3540_wire_157_7,
c3540_wire_157_8,
c3540_wire_157_9,
c3540_wire_157_10,
c3540_wire_157_11,
c3540_wire_157_12,
c3540_wire_157_13,
c3540_wire_157_14,
c3540_wire_157_15,
c3540_wire_161_0,
c3540_wire_161_1,
c3540_wire_161_2,
c3540_wire_161_3,
c3540_wire_161_4,
c3540_wire_161_5,
c3540_wire_161_6,
c3540_wire_161_7,
c3540_wire_161_8,
c3540_wire_161_9,
c3540_wire_161_10,
c3540_wire_161_11,
c3540_wire_161_12,
c3540_wire_161_13,
c3540_wire_161_14,
c3540_wire_161_15,
c3540_wire_163_0,
c3540_wire_163_1,
c3540_wire_163_2,
c3540_wire_163_3,
c3540_wire_163_4,
c3540_wire_163_5,
c3540_wire_163_6,
c3540_wire_163_7,
c3540_wire_181_0,
c3540_wire_181_1,
c3540_wire_181_2,
c3540_wire_181_3,
c3540_wire_181_4,
c3540_wire_181_5,
c3540_wire_181_6,
c3540_wire_181_7,
c3540_wire_181_8,
c3540_wire_181_9,
c3540_wire_181_10,
c3540_wire_181_11,
c3540_wire_181_12,
c3540_wire_181_13,
c3540_wire_192_0,
c3540_wire_192_1,
c3540_wire_198_0,
c3540_wire_198_1,
c3540_wire_200_0,
c3540_wire_200_1,
c3540_wire_200_2,
c3540_wire_200_3,
c3540_wire_215_0,
c3540_wire_215_1,
c3540_wire_215_2,
c3540_wire_215_3,
c3540_wire_224_0,
c3540_wire_224_1,
c3540_wire_224_2,
c3540_wire_224_3,
c3540_wire_224_4,
c3540_wire_224_5,
c3540_wire_224_6,
c3540_wire_224_7,
c3540_wire_224_8,
c3540_wire_224_9,
c3540_wire_224_10,
c3540_wire_224_11,
c3540_wire_224_12,
c3540_wire_224_13,
c3540_wire_224_14,
c3540_wire_224_15,
c3540_wire_242_0,
c3540_wire_242_1,
c3540_wire_242_2,
c3540_wire_242_3,
c3540_wire_242_4,
c3540_wire_242_5,
c3540_wire_242_6,
c3540_wire_242_7,
c3540_wire_242_8,
c3540_wire_242_9,
c3540_wire_242_10,
c3540_wire_242_11,
c3540_wire_242_12,
c3540_wire_242_13,
c3540_wire_242_14,
c3540_wire_242_15,
c3540_wire_298_0,
c3540_wire_298_1,
c3540_wire_45_0,
c3540_wire_45_1,
c3540_wire_45_2,
c3540_wire_45_3,
c3540_wire_327_0,
c3540_wire_327_1,
c3540_wire_327_2,
c3540_wire_350_0,
c3540_wire_350_1,
c3540_wire_350_2,
c3540_wire_352_0,
c3540_wire_352_1,
c3540_wire_352_2,
c3540_wire_367_0,
c3540_wire_367_1,
c3540_wire_367_2,
c3540_wire_73_0,
c3540_wire_73_1,
c3540_wire_73_2,
c3540_wire_73_3,
c3540_wire_73_4,
c3540_wire_388_0,
c3540_wire_388_1,
c3540_wire_388_2,
c3540_wire_403_0,
c3540_wire_403_1,
c3540_wire_75_0,
c3540_wire_75_1,
c3540_wire_75_2,
c3540_wire_75_3,
c3540_wire_75_4,
c3540_wire_417_0,
c3540_wire_417_1,
c3540_wire_417_2,
c3540_wire_69_0,
c3540_wire_69_1,
c3540_wire_69_2,
c3540_wire_69_3,
c3540_wire_69_4,
c3540_wire_450_0,
c3540_wire_450_1,
c3540_wire_450_2,
c3540_wire_450_3,
c3540_wire_450_4,
c3540_wire_454_0,
c3540_wire_454_1,
c3540_wire_454_2,
c3540_wire_454_3,
c3540_wire_454_4,
c3540_wire_493_0,
c3540_wire_493_1,
c3540_wire_493_2,
c3540_wire_79_0,
c3540_wire_79_1,
c3540_wire_79_2,
c3540_wire_79_3,
c3540_wire_79_4,
c3540_wire_455_0,
c3540_wire_455_1,
c3540_wire_455_2,
c3540_wire_455_3,
c3540_wire_455_4,
c3540_wire_525_0,
c3540_wire_525_1,
c3540_wire_525_2,
c3540_wire_71_0,
c3540_wire_71_1,
c3540_wire_71_2,
c3540_wire_71_3,
c3540_wire_71_4,
c3540_wire_456_0,
c3540_wire_456_1,
c3540_wire_456_2,
c3540_wire_456_3,
c3540_wire_456_4,
c3540_wire_566_0,
c3540_wire_566_1,
c3540_wire_566_2,
c3540_wire_566_3,
c3540_wire_221_0,
c3540_wire_221_1,
c3540_wire_221_2,
c3540_wire_221_3,
c3540_wire_297_0,
c3540_wire_297_1,
c3540_wire_297_2,
c3540_wire_297_3,
c3540_wire_297_4,
c3540_wire_325_0,
c3540_wire_325_1,
c3540_wire_325_2,
c3540_wire_325_3,
c3540_wire_325_4,
c3540_wire_325_5,
c3540_wire_325_6,
c3540_wire_325_7,
c3540_wire_325_8,
c3540_wire_325_9,
c3540_wire_325_10,
c3540_wire_325_11,
c3540_wire_325_12,
c3540_wire_325_13,
c3540_wire_325_14,
c3540_wire_325_15,
c3540_wire_325_16,
c3540_wire_325_17,
c3540_wire_325_18,
c3540_wire_32_0,
c3540_wire_32_1,
c3540_wire_32_2,
c3540_wire_32_3,
c3540_wire_32_4,
c3540_wire_32_5,
c3540_wire_32_6,
c3540_wire_32_7,
c3540_wire_32_8,
c3540_wire_32_9,
c3540_wire_32_10,
c3540_wire_32_11,
c3540_wire_32_12,
c3540_wire_32_13,
c3540_wire_32_14,
c3540_wire_32_15,
c3540_wire_32_16,
c3540_wire_32_17,
c3540_wire_32_18,
c3540_wire_32_19,
c3540_wire_32_20,
c3540_wire_32_21,
c3540_wire_32_22,
c3540_wire_349_0,
c3540_wire_349_1,
c3540_wire_349_2,
c3540_wire_349_3,
c3540_wire_349_4,
c3540_wire_349_5,
c3540_wire_596_0,
c3540_wire_596_1,
c3540_wire_138_0,
c3540_wire_138_1,
c3540_wire_313_0,
c3540_wire_313_1,
c3540_wire_313_2,
c3540_wire_313_3,
c3540_wire_313_4,
c3540_wire_313_5,
c3540_wire_313_6,
c3540_wire_313_7,
c3540_wire_572_0,
c3540_wire_572_1,
c3540_wire_572_2,
c3540_wire_572_3,
c3540_wire_572_4,
c3540_wire_572_5,
c3540_wire_572_6,
c3540_wire_572_7,
c3540_wire_572_8,
c3540_wire_694_0,
c3540_wire_694_1,
c3540_wire_47_0,
c3540_wire_47_1,
c3540_wire_47_2,
c3540_wire_47_3,
c3540_wire_715_0,
c3540_wire_715_1,
c3540_wire_77_0,
c3540_wire_77_1,
c3540_wire_77_2,
c3540_wire_77_3,
c3540_wire_77_4,
c3540_wire_178_0,
c3540_wire_178_1,
c3540_wire_178_2,
c3540_wire_178_3,
c3540_wire_178_4,
c3540_wire_178_5,
c3540_wire_178_6,
c3540_wire_178_7,
c3540_wire_178_8,
c3540_wire_178_9,
c3540_wire_178_10,
c3540_wire_178_11,
c3540_wire_178_12,
c3540_wire_178_13,
c3540_wire_178_14,
c3540_wire_178_15,
c3540_wire_178_16,
c3540_wire_733_0,
c3540_wire_733_1,
c3540_wire_733_2,
c3540_wire_738_0,
c3540_wire_738_1,
c3540_wire_738_2,
c3540_wire_732_0,
c3540_wire_732_1,
c3540_wire_732_2,
c3540_wire_732_3,
c3540_wire_732_4,
c3540_wire_732_5,
c3540_wire_732_6,
c3540_wire_732_7,
c3540_wire_150_0,
c3540_wire_150_1,
c3540_wire_150_2,
c3540_wire_150_3,
c3540_wire_150_4,
c3540_wire_150_5,
c3540_wire_150_6,
c3540_wire_150_7,
c3540_wire_150_8,
c3540_wire_150_9,
c3540_wire_150_10,
c3540_wire_150_11,
c3540_wire_150_12,
c3540_wire_150_13,
c3540_wire_150_14,
c3540_wire_150_15,
c3540_wire_150_16,
c3540_wire_150_17,
c3540_wire_150_18,
c3540_wire_150_19,
c3540_wire_150_20,
c3540_wire_150_21,
c3540_wire_150_22,
c3540_wire_741_0,
c3540_wire_741_1,
c3540_wire_741_2,
c3540_wire_741_3,
c3540_wire_741_4,
c3540_wire_741_5,
c3540_wire_597_0,
c3540_wire_597_1,
c3540_wire_597_2,
c3540_wire_742_0,
c3540_wire_742_1,
c3540_wire_742_2,
c3540_wire_742_3,
c3540_wire_743_0,
c3540_wire_743_1,
c3540_wire_743_2,
c3540_wire_743_3,
c3540_wire_82_0,
c3540_wire_82_1,
c3540_wire_82_2,
c3540_wire_82_3,
c3540_wire_82_4,
c3540_wire_83_0,
c3540_wire_83_1,
c3540_wire_83_2,
c3540_wire_83_3,
c3540_wire_83_4,
c3540_wire_83_5,
c3540_wire_84_0,
c3540_wire_84_1,
c3540_wire_84_2,
c3540_wire_84_3,
c3540_wire_782_0,
c3540_wire_782_1,
c3540_wire_782_2,
c3540_wire_782_3,
c3540_wire_159_0,
c3540_wire_159_1,
c3540_wire_149_0,
c3540_wire_149_1,
c3540_wire_149_2,
c3540_wire_149_3,
c3540_wire_149_4,
c3540_wire_149_5,
c3540_wire_149_6,
c3540_wire_149_7,
c3540_wire_149_8,
c3540_wire_149_9,
c3540_wire_149_10,
c3540_wire_149_11,
c3540_wire_149_12,
c3540_wire_740_0,
c3540_wire_740_1,
c3540_wire_740_2,
c3540_wire_85_0,
c3540_wire_85_1,
c3540_wire_85_2,
c3540_wire_85_3,
c3540_wire_85_4,
c3540_wire_85_5,
c3540_wire_158_0,
c3540_wire_158_1,
c3540_wire_151_0,
c3540_wire_151_1,
c3540_wire_151_2,
c3540_wire_151_3,
c3540_wire_151_4,
c3540_wire_151_5,
c3540_wire_151_6,
c3540_wire_151_7,
c3540_wire_151_8,
c3540_wire_151_9,
c3540_wire_151_10,
c3540_wire_151_11,
c3540_wire_151_12,
c3540_wire_151_13,
c3540_wire_805_0,
c3540_wire_805_1,
c3540_wire_807_0,
c3540_wire_807_1,
c3540_wire_807_2,
c3540_wire_815_0,
c3540_wire_815_1,
c3540_wire_815_2,
c3540_wire_815_3,
c3540_wire_815_4,
c3540_wire_815_5,
c3540_wire_815_6,
c3540_wire_815_7,
c3540_wire_815_8,
c3540_wire_815_9,
c3540_wire_827_0,
c3540_wire_827_1,
c3540_wire_827_2,
c3540_wire_827_3,
c3540_wire_827_4,
c3540_wire_827_5,
c3540_wire_827_6,
c3540_wire_41_0,
c3540_wire_41_1,
c3540_wire_41_2,
c3540_wire_41_3,
c3540_wire_41_4,
c3540_wire_41_5,
c3540_wire_836_0,
c3540_wire_836_1,
c3540_wire_799_0,
c3540_wire_799_1,
c3540_wire_799_2,
c3540_wire_799_3,
c3540_wire_799_4,
c3540_wire_799_5,
c3540_wire_799_6,
c3540_wire_799_7,
c3540_wire_799_8,
c3540_wire_799_9,
c3540_wire_800_0,
c3540_wire_800_1,
c3540_wire_800_2,
c3540_wire_800_3,
c3540_wire_800_4,
c3540_wire_800_5,
c3540_wire_800_6,
c3540_wire_800_7,
c3540_wire_800_8,
c3540_wire_855_0,
c3540_wire_855_1,
c3540_wire_855_2,
c3540_wire_785_0,
c3540_wire_785_1,
c3540_wire_785_2,
c3540_wire_785_3,
c3540_wire_785_4,
c3540_wire_785_5,
c3540_wire_785_6,
c3540_wire_864_0,
c3540_wire_864_1,
c3540_wire_864_2,
c3540_wire_864_3,
c3540_wire_864_4,
c3540_wire_864_5,
c3540_wire_864_6,
c3540_wire_864_7,
c3540_wire_904_0,
c3540_wire_904_1,
c3540_wire_904_2,
c3540_wire_904_3,
c3540_wire_904_4,
c3540_wire_909_0,
c3540_wire_909_1,
c3540_wire_909_2,
c3540_wire_909_3,
c3540_wire_909_4,
c3540_wire_916_0,
c3540_wire_916_1,
c3540_wire_917_0,
c3540_wire_917_1,
c3540_wire_935_0,
c3540_wire_935_1,
c3540_wire_935_2,
c3540_wire_935_3,
c3540_wire_938_0,
c3540_wire_938_1,
c3540_wire_942_0,
c3540_wire_942_1,
c3540_wire_942_2,
c3540_wire_942_3,
c3540_wire_940_0,
c3540_wire_940_1,
c3540_wire_333_0,
c3540_wire_333_1,
c3540_wire_943_0,
c3540_wire_943_1,
c3540_wire_943_2,
c3540_wire_943_3,
c3540_wire_946_0,
c3540_wire_946_1,
c3540_wire_946_2,
c3540_wire_952_0,
c3540_wire_952_1,
c3540_wire_913_0,
c3540_wire_913_1,
c3540_wire_913_2,
c3540_wire_913_3,
c3540_wire_837_0,
c3540_wire_837_1,
c3540_wire_958_0,
c3540_wire_958_1,
c3540_wire_33_0,
c3540_wire_33_1,
c3540_wire_33_2,
c3540_wire_33_3,
c3540_wire_33_4,
c3540_wire_33_5,
c3540_wire_33_6,
c3540_wire_33_7,
c3540_wire_33_8,
c3540_wire_33_9,
c3540_wire_33_10,
c3540_wire_33_11,
c3540_wire_33_12,
c3540_wire_33_13,
c3540_wire_33_14,
c3540_wire_33_15,
c3540_wire_33_16,
c3540_wire_33_17,
c3540_wire_33_18,
c3540_wire_33_19,
c3540_wire_33_20,
c3540_wire_33_21,
c3540_wire_33_22,
c3540_wire_33_23,
c3540_wire_33_24,
c3540_wire_33_25,
c3540_wire_33_26,
c3540_wire_33_27,
c3540_wire_33_28,
c3540_wire_33_29,
c3540_wire_33_30,
c3540_wire_33_31,
c3540_wire_33_32,
c3540_wire_33_33,
c3540_wire_33_34,
c3540_wire_33_35,
c3540_wire_33_36,
c3540_wire_33_37,
c3540_wire_33_38,
c3540_wire_33_39,
c3540_wire_9_0,
c3540_wire_9_1,
c3540_wire_9_2,
c3540_wire_9_3,
c3540_wire_9_4,
c3540_wire_9_5,
c3540_wire_973_0,
c3540_wire_973_1,
c3540_wire_973_2,
c3540_wire_973_3,
c3540_wire_10_0,
c3540_wire_10_1,
c3540_wire_10_2,
c3540_wire_10_3,
c3540_wire_10_4,
c3540_wire_10_5,
c3540_wire_1019_0,
c3540_wire_1019_1,
c3540_wire_1019_2,
c3540_wire_1019_3,
c3540_wire_1019_4,
c3540_wire_1023_0,
c3540_wire_1023_1,
c3540_wire_1023_2,
c3540_wire_1023_3,
c3540_wire_1028_0,
c3540_wire_1028_1,
c3540_wire_1028_2,
c3540_wire_1028_3,
c3540_wire_1030_0,
c3540_wire_1030_1,
c3540_wire_824_0,
c3540_wire_824_1,
c3540_wire_824_2,
c3540_wire_824_3,
c3540_wire_824_4,
c3540_wire_1045_0,
c3540_wire_1045_1,
c3540_wire_1045_2,
c3540_wire_1045_3,
c3540_wire_401_0,
c3540_wire_401_1,
c3540_wire_401_2,
c3540_wire_401_3,
c3540_wire_401_4,
c3540_wire_401_5,
c3540_wire_401_6,
c3540_wire_401_7,
c3540_wire_976_0,
c3540_wire_976_1,
c3540_wire_976_2,
c3540_wire_976_3,
c3540_wire_976_4,
c3540_wire_1104_0,
c3540_wire_1104_1,
c3540_wire_1104_2,
c3540_wire_1104_3,
c3540_wire_1104_4,
c3540_wire_1104_5,
c3540_wire_1104_6,
c3540_wire_1122_0,
c3540_wire_1122_1,
c3540_wire_1122_2,
c3540_wire_1122_3,
c3540_wire_1122_4,
c3540_wire_1159_0,
c3540_wire_1159_1,
c3540_wire_1159_2,
c3540_wire_1159_3,
c3540_wire_1159_4,
c3540_wire_1159_5,
c3540_wire_1159_6,
c3540_wire_430_0,
c3540_wire_430_1,
c3540_wire_430_2,
c3540_wire_430_3,
c3540_wire_430_4,
c3540_wire_430_5,
c3540_wire_430_6,
c3540_wire_430_7,
c3540_wire_1167_0,
c3540_wire_1167_1,
c3540_wire_1167_2,
c3540_wire_1167_3,
c3540_wire_1167_4,
c3540_wire_1167_5,
c3540_wire_1173_0,
c3540_wire_1173_1,
c3540_wire_1173_2,
c3540_wire_1173_3,
c3540_wire_1180_0,
c3540_wire_1180_1,
c3540_wire_1180_2,
c3540_wire_1180_3,
c3540_wire_1180_4,
c3540_wire_1180_5,
c3540_wire_1186_0,
c3540_wire_1186_1,
c3540_wire_28_0,
c3540_wire_28_1,
c3540_wire_28_2,
c3540_wire_28_3,
c3540_wire_28_4,
c3540_wire_28_5,
c3540_wire_28_6,
c3540_wire_1193_0,
c3540_wire_1193_1,
c3540_wire_1195_0,
c3540_wire_1195_1,
c3540_wire_1195_2,
c3540_wire_1195_3,
c3540_wire_1196_0,
c3540_wire_1196_1,
c3540_wire_1200_0,
c3540_wire_1200_1,
c3540_wire_1200_2,
c3540_wire_111_0,
c3540_wire_111_1,
c3540_wire_111_2,
c3540_wire_111_3,
c3540_wire_111_4,
c3540_wire_111_5,
c3540_wire_111_6,
c3540_wire_115_0,
c3540_wire_115_1,
c3540_wire_115_2,
c3540_wire_115_3,
c3540_wire_115_4,
c3540_wire_115_5,
c3540_wire_116_0,
c3540_wire_116_1,
c3540_wire_116_2,
c3540_wire_116_3,
c3540_wire_340_0,
c3540_wire_340_1,
c3540_wire_340_2,
c3540_wire_340_3,
c3540_wire_340_4,
c3540_wire_340_5,
c3540_wire_340_6,
c3540_wire_340_7,
c3540_wire_483_0,
c3540_wire_483_1,
c3540_wire_483_2,
c3540_wire_483_3,
c3540_wire_483_4,
c3540_wire_483_5,
c3540_wire_483_6,
c3540_wire_483_7,
c3540_wire_483_8,
c3540_wire_326_0,
c3540_wire_326_1,
c3540_wire_326_2,
c3540_wire_326_3,
c3540_wire_60_0,
c3540_wire_60_1,
c3540_wire_60_2,
c3540_wire_60_3,
c3540_wire_60_4,
c3540_wire_60_5,
c3540_wire_60_6,
c3540_wire_60_7,
c3540_wire_60_8,
c3540_wire_60_9,
c3540_wire_60_10,
c3540_wire_60_11,
c3540_wire_60_12,
c3540_wire_60_13,
c3540_wire_60_14,
c3540_wire_60_15,
c3540_wire_60_16,
c3540_wire_60_17,
c3540_wire_60_18,
c3540_wire_60_19,
c3540_wire_60_20,
c3540_wire_60_21,
c3540_wire_60_22,
c3540_wire_60_23,
c3540_wire_60_24,
c3540_wire_60_25,
c3540_wire_60_26,
c3540_wire_60_27,
c3540_wire_60_28,
c3540_wire_60_29,
c3540_wire_60_30,
c3540_wire_60_31,
c3540_wire_60_32,
c3540_wire_60_33,
c3540_wire_60_34,
c3540_wire_60_35,
c3540_wire_60_36,
c3540_wire_60_37,
c3540_wire_60_38,
c3540_wire_60_39,
c3540_wire_60_40,
c3540_wire_60_41,
c3540_wire_60_42,
c3540_wire_60_43,
c3540_wire_60_44,
c3540_wire_60_45,
c3540_wire_60_46,
c3540_wire_60_47,
c3540_wire_60_48,
c3540_wire_60_49,
c3540_wire_60_50,
c3540_wire_60_51,
c3540_wire_60_52,
c3540_wire_60_53,
c3540_wire_60_54,
c3540_wire_516_0,
c3540_wire_516_1,
c3540_wire_516_2,
c3540_wire_516_3,
c3540_wire_516_4,
c3540_wire_516_5,
c3540_wire_516_6,
c3540_wire_549_0,
c3540_wire_549_1,
c3540_wire_549_2,
c3540_wire_549_3,
c3540_wire_549_4,
c3540_wire_549_5,
c3540_wire_549_6,
c3540_wire_685_0,
c3540_wire_685_1,
c3540_wire_685_2,
c3540_wire_685_3,
c3540_wire_685_4,
c3540_wire_1002_0,
c3540_wire_1002_1,
c3540_wire_1002_2,
c3540_wire_1002_3,
c3540_wire_994_0,
c3540_wire_994_1,
c3540_wire_994_2,
c3540_wire_997_0,
c3540_wire_997_1,
c3540_wire_832_0,
c3540_wire_832_1,
c3540_wire_832_2,
c3540_wire_832_3,
c3540_wire_832_4,
c3540_wire_832_5,
c3540_wire_832_6,
c3540_wire_832_7,
c3540_wire_832_8,
c3540_wire_832_9,
c3540_wire_832_10,
c3540_wire_832_11,
c3540_wire_832_12,
c3540_wire_832_13,
c3540_wire_832_14,
c3540_wire_42_0,
c3540_wire_42_1,
c3540_wire_344_0,
c3540_wire_344_1,
c3540_wire_344_2,
c3540_wire_344_3,
c3540_wire_344_4,
c3540_wire_344_5,
c3540_wire_344_6,
c3540_wire_344_7,
c3540_wire_449_0,
c3540_wire_449_1,
c3540_wire_449_2,
c3540_wire_449_3,
c3540_wire_38_0,
c3540_wire_38_1,
c3540_wire_38_2,
c3540_wire_38_3,
c3540_wire_38_4,
c3540_wire_38_5,
c3540_wire_38_6,
c3540_wire_38_7,
c3540_wire_38_8,
c3540_wire_38_9,
c3540_wire_38_10,
c3540_wire_38_11,
c3540_wire_38_12,
c3540_wire_38_13,
c3540_wire_38_14,
c3540_wire_38_15,
c3540_wire_38_16,
c3540_wire_469_0,
c3540_wire_469_1,
c3540_wire_469_2,
c3540_wire_469_3,
c3540_wire_469_4,
c3540_wire_469_5,
c3540_wire_469_6,
c3540_wire_469_7,
c3540_wire_469_8,
c3540_wire_469_9,
c3540_wire_469_10,
c3540_wire_469_11,
c3540_wire_1049_0,
c3540_wire_1049_1,
c3540_wire_1049_2,
c3540_wire_1049_3,
c3540_wire_1049_4,
c3540_wire_18_0,
c3540_wire_18_1,
c3540_wire_18_2,
c3540_wire_18_3,
c3540_wire_18_4,
c3540_wire_18_5,
c3540_wire_18_6,
c3540_wire_18_7,
c3540_wire_18_8,
c3540_wire_18_9,
c3540_wire_18_10,
c3540_wire_18_11,
c3540_wire_18_12,
c3540_wire_18_13,
c3540_wire_18_14,
c3540_wire_18_15,
c3540_wire_18_16,
c3540_wire_18_17,
c3540_wire_18_18,
c3540_wire_309_0,
c3540_wire_309_1,
c3540_wire_341_0,
c3540_wire_341_1,
c3540_wire_341_2,
c3540_wire_341_3,
c3540_wire_341_4,
c3540_wire_341_5,
c3540_wire_341_6,
c3540_wire_341_7,
c3540_wire_492_0,
c3540_wire_492_1,
c3540_wire_492_2,
c3540_wire_120_0,
c3540_wire_120_1,
c3540_wire_120_2,
c3540_wire_120_3,
c3540_wire_120_4,
c3540_wire_120_5,
c3540_wire_120_6,
c3540_wire_120_7,
c3540_wire_120_8,
c3540_wire_120_9,
c3540_wire_120_10,
c3540_wire_120_11,
c3540_wire_120_12,
c3540_wire_120_13,
c3540_wire_120_14,
c3540_wire_120_15,
c3540_wire_120_16,
c3540_wire_120_17,
c3540_wire_120_18,
c3540_wire_318_0,
c3540_wire_318_1,
c3540_wire_318_2,
c3540_wire_318_3,
c3540_wire_318_4,
c3540_wire_318_5,
c3540_wire_318_6,
c3540_wire_318_7,
c3540_wire_318_8,
c3540_wire_318_9,
c3540_wire_318_10,
c3540_wire_318_11,
c3540_wire_318_12,
c3540_wire_318_13,
c3540_wire_318_14,
c3540_wire_318_15,
c3540_wire_121_0,
c3540_wire_121_1,
c3540_wire_121_2,
c3540_wire_121_3,
c3540_wire_121_4,
c3540_wire_121_5,
c3540_wire_121_6,
c3540_wire_121_7,
c3540_wire_121_8,
c3540_wire_121_9,
c3540_wire_121_10,
c3540_wire_121_11,
c3540_wire_121_12,
c3540_wire_121_13,
c3540_wire_121_14,
c3540_wire_121_15,
c3540_wire_121_16,
c3540_wire_121_17,
c3540_wire_121_18,
c3540_wire_121_19,
c3540_wire_121_20,
c3540_wire_121_21,
c3540_wire_121_22,
c3540_wire_1009_0,
c3540_wire_1009_1,
c3540_wire_1009_2,
c3540_wire_1009_3,
c3540_wire_1009_4,
c3540_wire_1009_5,
c3540_wire_1009_6,
c3540_wire_1009_7,
c3540_wire_346_0,
c3540_wire_346_1,
c3540_wire_346_2,
c3540_wire_346_3,
c3540_wire_346_4,
c3540_wire_346_5,
c3540_wire_346_6,
c3540_wire_346_7,
G1_net_0,
G2_net_0,
G3_net_0,
G4_net_0,
G5_net_0,
G6_net_0,
G7_net_0,
G8_net_0,
G9_net_0,
G10_net_0,
G11_net_0,
G12_net_0,
G13_net_0,
G14_net_0,
G15_net_0,
G16_net_0,
G17_net_0,
G18_net_0,
G19_net_0,
G20_net_0,
G21_net_0,
G22_net_0,
G23_net_0,
G24_net_0,
G25_net_0,
G26_net_0,
G27_net_0,
G28_net_0,
G29_net_0,
G30_net_0,
G31_net_0,
G32_net_0,
G33_net_0,
G34_net_0,
G35_net_0,
G36_net_0,
G37_net_0,
G38_net_0,
G39_net_0,
G40_net_0,
G41_net_0,
G42_net_0,
G43_net_0,
G44_net_0,
G45_net_0,
G46_net_0,
G47_net_0,
G48_net_0,
G49_net_0,
G50_net_0,
G3519_net_0,
G3520_net_0,
G3521_net_0,
G3522_net_0,
G3523_net_0,
G3524_net_0,
G3525_net_0,
G3526_net_0,
G3527_net_0,
G3528_net_0,
G3529_net_0,
G3530_net_0,
G3531_net_0,
G3532_net_0,
G3533_net_0,
G3534_net_0,
G3535_net_0,
G3536_net_0,
G3537_net_0,
G3538_net_0,
G3539_net_0,
G3540_net_0;

pin #(50) pin_0 ({G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G50}, {G1_net_0, G2_net_0, G3_net_0, G4_net_0, G5_net_0, G6_net_0, G7_net_0, G8_net_0, G9_net_0, G10_net_0, G11_net_0, G12_net_0, G13_net_0, G14_net_0, G15_net_0, G16_net_0, G17_net_0, G18_net_0, G19_net_0, G20_net_0, G21_net_0, G22_net_0, G23_net_0, G24_net_0, G25_net_0, G26_net_0, G27_net_0, G28_net_0, G29_net_0, G30_net_0, G31_net_0, G32_net_0, G33_net_0, G34_net_0, G35_net_0, G36_net_0, G37_net_0, G38_net_0, G39_net_0, G40_net_0, G41_net_0, G42_net_0, G43_net_0, G44_net_0, G45_net_0, G46_net_0, G47_net_0, G48_net_0, G49_net_0, G50_net_0});

pout #(22) pout_0 ({G3519_net_0, G3520_net_0, G3521_net_0, G3522_net_0, G3523_net_0, G3524_net_0, G3525_net_0, G3526_net_0, G3527_net_0, G3528_net_0, G3529_net_0, G3530_net_0, G3531_net_0, G3532_net_0, G3533_net_0, G3534_net_0, G3535_net_0, G3536_net_0, G3537_net_0, G3538_net_0, G3539_net_0, G3540_net_0}, {G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540});

fanout_n #(28, 0, 0) FANOUT_1 (c3540_wire_1, {c3540_wire_1_0, c3540_wire_1_1, c3540_wire_1_2, c3540_wire_1_3, c3540_wire_1_4, c3540_wire_1_5, c3540_wire_1_6, c3540_wire_1_7, c3540_wire_1_8, c3540_wire_1_9, c3540_wire_1_10, c3540_wire_1_11, c3540_wire_1_12, c3540_wire_1_13, c3540_wire_1_14, c3540_wire_1_15, c3540_wire_1_16, c3540_wire_1_17, c3540_wire_1_18, c3540_wire_1_19, c3540_wire_1_20, c3540_wire_1_21, c3540_wire_1_22, c3540_wire_1_23, c3540_wire_1_24, c3540_wire_1_25, c3540_wire_1_26, c3540_wire_1_27});
fanout_n #(17, 0, 0) FANOUT_2 (c3540_wire_2, {c3540_wire_2_0, c3540_wire_2_1, c3540_wire_2_2, c3540_wire_2_3, c3540_wire_2_4, c3540_wire_2_5, c3540_wire_2_6, c3540_wire_2_7, c3540_wire_2_8, c3540_wire_2_9, c3540_wire_2_10, c3540_wire_2_11, c3540_wire_2_12, c3540_wire_2_13, c3540_wire_2_14, c3540_wire_2_15, c3540_wire_2_16});
fanout_n #(2, 0, 0) FANOUT_3 (c3540_wire_11, {c3540_wire_11_0, c3540_wire_11_1});
fanout_n #(2, 0, 0) FANOUT_4 (c3540_wire_30, {c3540_wire_30_0, c3540_wire_30_1});
fanout_n #(9, 0, 0) FANOUT_5 (c3540_wire_35, {c3540_wire_35_0, c3540_wire_35_1, c3540_wire_35_2, c3540_wire_35_3, c3540_wire_35_4, c3540_wire_35_5, c3540_wire_35_6, c3540_wire_35_7, c3540_wire_35_8});
fanout_n #(6, 0, 0) FANOUT_6 (c3540_wire_39, {c3540_wire_39_0, c3540_wire_39_1, c3540_wire_39_2, c3540_wire_39_3, c3540_wire_39_4, c3540_wire_39_5});
fanout_n #(23, 0, 0) FANOUT_7 (c3540_wire_40, {c3540_wire_40_0, c3540_wire_40_1, c3540_wire_40_2, c3540_wire_40_3, c3540_wire_40_4, c3540_wire_40_5, c3540_wire_40_6, c3540_wire_40_7, c3540_wire_40_8, c3540_wire_40_9, c3540_wire_40_10, c3540_wire_40_11, c3540_wire_40_12, c3540_wire_40_13, c3540_wire_40_14, c3540_wire_40_15, c3540_wire_40_16, c3540_wire_40_17, c3540_wire_40_18, c3540_wire_40_19, c3540_wire_40_20, c3540_wire_40_21, c3540_wire_40_22});
fanout_n #(16, 0, 0) FANOUT_8 (c3540_wire_5, {c3540_wire_5_0, c3540_wire_5_1, c3540_wire_5_2, c3540_wire_5_3, c3540_wire_5_4, c3540_wire_5_5, c3540_wire_5_6, c3540_wire_5_7, c3540_wire_5_8, c3540_wire_5_9, c3540_wire_5_10, c3540_wire_5_11, c3540_wire_5_12, c3540_wire_5_13, c3540_wire_5_14, c3540_wire_5_15});
fanout_n #(3, 0, 0) FANOUT_9 (c3540_wire_93, {c3540_wire_93_0, c3540_wire_93_1, c3540_wire_93_2});
fanout_n #(17, 0, 0) FANOUT_10 (c3540_wire_99, {c3540_wire_99_0, c3540_wire_99_1, c3540_wire_99_2, c3540_wire_99_3, c3540_wire_99_4, c3540_wire_99_5, c3540_wire_99_6, c3540_wire_99_7, c3540_wire_99_8, c3540_wire_99_9, c3540_wire_99_10, c3540_wire_99_11, c3540_wire_99_12, c3540_wire_99_13, c3540_wire_99_14, c3540_wire_99_15, c3540_wire_99_16});
fanout_n #(2, 0, 0) FANOUT_11 (c3540_wire_112, {c3540_wire_112_0, c3540_wire_112_1});
fanout_n #(2, 0, 0) FANOUT_12 (c3540_wire_117, {c3540_wire_117_0, c3540_wire_117_1});
fanout_n #(2, 0, 0) FANOUT_13 (c3540_wire_119, {c3540_wire_119_0, c3540_wire_119_1});
fanout_n #(2, 0, 0) FANOUT_14 (c3540_wire_125, {c3540_wire_125_0, c3540_wire_125_1});
fanout_n #(16, 0, 0) FANOUT_15 (c3540_wire_123, {c3540_wire_123_0, c3540_wire_123_1, c3540_wire_123_2, c3540_wire_123_3, c3540_wire_123_4, c3540_wire_123_5, c3540_wire_123_6, c3540_wire_123_7, c3540_wire_123_8, c3540_wire_123_9, c3540_wire_123_10, c3540_wire_123_11, c3540_wire_123_12, c3540_wire_123_13, c3540_wire_123_14, c3540_wire_123_15});
fanout_n #(8, 0, 0) FANOUT_16 (c3540_wire_153, {c3540_wire_153_0, c3540_wire_153_1, c3540_wire_153_2, c3540_wire_153_3, c3540_wire_153_4, c3540_wire_153_5, c3540_wire_153_6, c3540_wire_153_7});
fanout_n #(16, 0, 0) FANOUT_17 (c3540_wire_155, {c3540_wire_155_0, c3540_wire_155_1, c3540_wire_155_2, c3540_wire_155_3, c3540_wire_155_4, c3540_wire_155_5, c3540_wire_155_6, c3540_wire_155_7, c3540_wire_155_8, c3540_wire_155_9, c3540_wire_155_10, c3540_wire_155_11, c3540_wire_155_12, c3540_wire_155_13, c3540_wire_155_14, c3540_wire_155_15});
fanout_n #(16, 0, 0) FANOUT_18 (c3540_wire_157, {c3540_wire_157_0, c3540_wire_157_1, c3540_wire_157_2, c3540_wire_157_3, c3540_wire_157_4, c3540_wire_157_5, c3540_wire_157_6, c3540_wire_157_7, c3540_wire_157_8, c3540_wire_157_9, c3540_wire_157_10, c3540_wire_157_11, c3540_wire_157_12, c3540_wire_157_13, c3540_wire_157_14, c3540_wire_157_15});
fanout_n #(16, 0, 0) FANOUT_19 (c3540_wire_161, {c3540_wire_161_0, c3540_wire_161_1, c3540_wire_161_2, c3540_wire_161_3, c3540_wire_161_4, c3540_wire_161_5, c3540_wire_161_6, c3540_wire_161_7, c3540_wire_161_8, c3540_wire_161_9, c3540_wire_161_10, c3540_wire_161_11, c3540_wire_161_12, c3540_wire_161_13, c3540_wire_161_14, c3540_wire_161_15});
fanout_n #(8, 0, 0) FANOUT_20 (c3540_wire_163, {c3540_wire_163_0, c3540_wire_163_1, c3540_wire_163_2, c3540_wire_163_3, c3540_wire_163_4, c3540_wire_163_5, c3540_wire_163_6, c3540_wire_163_7});
fanout_n #(14, 0, 0) FANOUT_21 (c3540_wire_181, {c3540_wire_181_0, c3540_wire_181_1, c3540_wire_181_2, c3540_wire_181_3, c3540_wire_181_4, c3540_wire_181_5, c3540_wire_181_6, c3540_wire_181_7, c3540_wire_181_8, c3540_wire_181_9, c3540_wire_181_10, c3540_wire_181_11, c3540_wire_181_12, c3540_wire_181_13});
fanout_n #(2, 0, 0) FANOUT_22 (c3540_wire_192, {c3540_wire_192_0, c3540_wire_192_1});
fanout_n #(2, 0, 0) FANOUT_23 (c3540_wire_198, {c3540_wire_198_0, c3540_wire_198_1});
fanout_n #(4, 0, 0) FANOUT_24 (c3540_wire_200, {c3540_wire_200_0, c3540_wire_200_1, c3540_wire_200_2, c3540_wire_200_3});
fanout_n #(4, 0, 0) FANOUT_25 (c3540_wire_215, {c3540_wire_215_0, c3540_wire_215_1, c3540_wire_215_2, c3540_wire_215_3});
fanout_n #(16, 0, 0) FANOUT_26 (c3540_wire_224, {c3540_wire_224_0, c3540_wire_224_1, c3540_wire_224_2, c3540_wire_224_3, c3540_wire_224_4, c3540_wire_224_5, c3540_wire_224_6, c3540_wire_224_7, c3540_wire_224_8, c3540_wire_224_9, c3540_wire_224_10, c3540_wire_224_11, c3540_wire_224_12, c3540_wire_224_13, c3540_wire_224_14, c3540_wire_224_15});
fanout_n #(16, 0, 0) FANOUT_27 (c3540_wire_242, {c3540_wire_242_0, c3540_wire_242_1, c3540_wire_242_2, c3540_wire_242_3, c3540_wire_242_4, c3540_wire_242_5, c3540_wire_242_6, c3540_wire_242_7, c3540_wire_242_8, c3540_wire_242_9, c3540_wire_242_10, c3540_wire_242_11, c3540_wire_242_12, c3540_wire_242_13, c3540_wire_242_14, c3540_wire_242_15});
fanout_n #(2, 0, 0) FANOUT_28 (c3540_wire_298, {c3540_wire_298_0, c3540_wire_298_1});
fanout_n #(4, 0, 0) FANOUT_29 (c3540_wire_45, {c3540_wire_45_0, c3540_wire_45_1, c3540_wire_45_2, c3540_wire_45_3});
fanout_n #(3, 0, 0) FANOUT_30 (c3540_wire_327, {c3540_wire_327_0, c3540_wire_327_1, c3540_wire_327_2});
fanout_n #(3, 0, 0) FANOUT_31 (c3540_wire_350, {c3540_wire_350_0, c3540_wire_350_1, c3540_wire_350_2});
fanout_n #(3, 0, 0) FANOUT_32 (c3540_wire_352, {c3540_wire_352_0, c3540_wire_352_1, c3540_wire_352_2});
fanout_n #(3, 0, 0) FANOUT_33 (c3540_wire_367, {c3540_wire_367_0, c3540_wire_367_1, c3540_wire_367_2});
fanout_n #(5, 0, 0) FANOUT_34 (c3540_wire_73, {c3540_wire_73_0, c3540_wire_73_1, c3540_wire_73_2, c3540_wire_73_3, c3540_wire_73_4});
fanout_n #(3, 0, 0) FANOUT_35 (c3540_wire_388, {c3540_wire_388_0, c3540_wire_388_1, c3540_wire_388_2});
fanout_n #(2, 0, 0) FANOUT_36 (c3540_wire_403, {c3540_wire_403_0, c3540_wire_403_1});
fanout_n #(5, 0, 0) FANOUT_37 (c3540_wire_75, {c3540_wire_75_0, c3540_wire_75_1, c3540_wire_75_2, c3540_wire_75_3, c3540_wire_75_4});
fanout_n #(3, 0, 0) FANOUT_38 (c3540_wire_417, {c3540_wire_417_0, c3540_wire_417_1, c3540_wire_417_2});
fanout_n #(5, 0, 0) FANOUT_39 (c3540_wire_69, {c3540_wire_69_0, c3540_wire_69_1, c3540_wire_69_2, c3540_wire_69_3, c3540_wire_69_4});
fanout_n #(5, 0, 0) FANOUT_40 (c3540_wire_450, {c3540_wire_450_0, c3540_wire_450_1, c3540_wire_450_2, c3540_wire_450_3, c3540_wire_450_4});
fanout_n #(5, 0, 0) FANOUT_41 (c3540_wire_454, {c3540_wire_454_0, c3540_wire_454_1, c3540_wire_454_2, c3540_wire_454_3, c3540_wire_454_4});
fanout_n #(3, 0, 0) FANOUT_42 (c3540_wire_493, {c3540_wire_493_0, c3540_wire_493_1, c3540_wire_493_2});
fanout_n #(5, 0, 0) FANOUT_43 (c3540_wire_79, {c3540_wire_79_0, c3540_wire_79_1, c3540_wire_79_2, c3540_wire_79_3, c3540_wire_79_4});
fanout_n #(5, 0, 0) FANOUT_44 (c3540_wire_455, {c3540_wire_455_0, c3540_wire_455_1, c3540_wire_455_2, c3540_wire_455_3, c3540_wire_455_4});
fanout_n #(3, 0, 0) FANOUT_45 (c3540_wire_525, {c3540_wire_525_0, c3540_wire_525_1, c3540_wire_525_2});
fanout_n #(5, 0, 0) FANOUT_46 (c3540_wire_71, {c3540_wire_71_0, c3540_wire_71_1, c3540_wire_71_2, c3540_wire_71_3, c3540_wire_71_4});
fanout_n #(5, 0, 0) FANOUT_47 (c3540_wire_456, {c3540_wire_456_0, c3540_wire_456_1, c3540_wire_456_2, c3540_wire_456_3, c3540_wire_456_4});
fanout_n #(4, 0, 0) FANOUT_48 (c3540_wire_566, {c3540_wire_566_0, c3540_wire_566_1, c3540_wire_566_2, c3540_wire_566_3});
fanout_n #(4, 0, 0) FANOUT_49 (c3540_wire_221, {c3540_wire_221_0, c3540_wire_221_1, c3540_wire_221_2, c3540_wire_221_3});
fanout_n #(5, 0, 0) FANOUT_50 (c3540_wire_297, {c3540_wire_297_0, c3540_wire_297_1, c3540_wire_297_2, c3540_wire_297_3, c3540_wire_297_4});
fanout_n #(19, 0, 0) FANOUT_51 (c3540_wire_325, {c3540_wire_325_0, c3540_wire_325_1, c3540_wire_325_2, c3540_wire_325_3, c3540_wire_325_4, c3540_wire_325_5, c3540_wire_325_6, c3540_wire_325_7, c3540_wire_325_8, c3540_wire_325_9, c3540_wire_325_10, c3540_wire_325_11, c3540_wire_325_12, c3540_wire_325_13, c3540_wire_325_14, c3540_wire_325_15, c3540_wire_325_16, c3540_wire_325_17, c3540_wire_325_18});
fanout_n #(23, 0, 0) FANOUT_52 (c3540_wire_32, {c3540_wire_32_0, c3540_wire_32_1, c3540_wire_32_2, c3540_wire_32_3, c3540_wire_32_4, c3540_wire_32_5, c3540_wire_32_6, c3540_wire_32_7, c3540_wire_32_8, c3540_wire_32_9, c3540_wire_32_10, c3540_wire_32_11, c3540_wire_32_12, c3540_wire_32_13, c3540_wire_32_14, c3540_wire_32_15, c3540_wire_32_16, c3540_wire_32_17, c3540_wire_32_18, c3540_wire_32_19, c3540_wire_32_20, c3540_wire_32_21, c3540_wire_32_22});
fanout_n #(6, 0, 0) FANOUT_53 (c3540_wire_349, {c3540_wire_349_0, c3540_wire_349_1, c3540_wire_349_2, c3540_wire_349_3, c3540_wire_349_4, c3540_wire_349_5});
fanout_n #(2, 0, 0) FANOUT_54 (c3540_wire_596, {c3540_wire_596_0, c3540_wire_596_1});
fanout_n #(2, 0, 0) FANOUT_55 (c3540_wire_138, {c3540_wire_138_0, c3540_wire_138_1});
fanout_n #(8, 0, 0) FANOUT_56 (c3540_wire_313, {c3540_wire_313_0, c3540_wire_313_1, c3540_wire_313_2, c3540_wire_313_3, c3540_wire_313_4, c3540_wire_313_5, c3540_wire_313_6, c3540_wire_313_7});
fanout_n #(9, 0, 0) FANOUT_57 (c3540_wire_572, {c3540_wire_572_0, c3540_wire_572_1, c3540_wire_572_2, c3540_wire_572_3, c3540_wire_572_4, c3540_wire_572_5, c3540_wire_572_6, c3540_wire_572_7, c3540_wire_572_8});
fanout_n #(2, 0, 0) FANOUT_58 (c3540_wire_694, {c3540_wire_694_0, c3540_wire_694_1});
fanout_n #(4, 0, 0) FANOUT_59 (c3540_wire_47, {c3540_wire_47_0, c3540_wire_47_1, c3540_wire_47_2, c3540_wire_47_3});
fanout_n #(2, 0, 0) FANOUT_60 (c3540_wire_715, {c3540_wire_715_0, c3540_wire_715_1});
fanout_n #(5, 0, 0) FANOUT_61 (c3540_wire_77, {c3540_wire_77_0, c3540_wire_77_1, c3540_wire_77_2, c3540_wire_77_3, c3540_wire_77_4});
fanout_n #(17, 0, 0) FANOUT_62 (c3540_wire_178, {c3540_wire_178_0, c3540_wire_178_1, c3540_wire_178_2, c3540_wire_178_3, c3540_wire_178_4, c3540_wire_178_5, c3540_wire_178_6, c3540_wire_178_7, c3540_wire_178_8, c3540_wire_178_9, c3540_wire_178_10, c3540_wire_178_11, c3540_wire_178_12, c3540_wire_178_13, c3540_wire_178_14, c3540_wire_178_15, c3540_wire_178_16});
fanout_n #(3, 0, 0) FANOUT_63 (c3540_wire_733, {c3540_wire_733_0, c3540_wire_733_1, c3540_wire_733_2});
fanout_n #(3, 0, 0) FANOUT_64 (c3540_wire_738, {c3540_wire_738_0, c3540_wire_738_1, c3540_wire_738_2});
fanout_n #(8, 0, 0) FANOUT_65 (c3540_wire_732, {c3540_wire_732_0, c3540_wire_732_1, c3540_wire_732_2, c3540_wire_732_3, c3540_wire_732_4, c3540_wire_732_5, c3540_wire_732_6, c3540_wire_732_7});
fanout_n #(23, 0, 0) FANOUT_66 (c3540_wire_150, {c3540_wire_150_0, c3540_wire_150_1, c3540_wire_150_2, c3540_wire_150_3, c3540_wire_150_4, c3540_wire_150_5, c3540_wire_150_6, c3540_wire_150_7, c3540_wire_150_8, c3540_wire_150_9, c3540_wire_150_10, c3540_wire_150_11, c3540_wire_150_12, c3540_wire_150_13, c3540_wire_150_14, c3540_wire_150_15, c3540_wire_150_16, c3540_wire_150_17, c3540_wire_150_18, c3540_wire_150_19, c3540_wire_150_20, c3540_wire_150_21, c3540_wire_150_22});
fanout_n #(6, 0, 0) FANOUT_67 (c3540_wire_741, {c3540_wire_741_0, c3540_wire_741_1, c3540_wire_741_2, c3540_wire_741_3, c3540_wire_741_4, c3540_wire_741_5});
fanout_n #(3, 0, 0) FANOUT_68 (c3540_wire_597, {c3540_wire_597_0, c3540_wire_597_1, c3540_wire_597_2});
fanout_n #(4, 0, 0) FANOUT_69 (c3540_wire_742, {c3540_wire_742_0, c3540_wire_742_1, c3540_wire_742_2, c3540_wire_742_3});
fanout_n #(4, 0, 0) FANOUT_70 (c3540_wire_743, {c3540_wire_743_0, c3540_wire_743_1, c3540_wire_743_2, c3540_wire_743_3});
fanout_n #(5, 0, 0) FANOUT_71 (c3540_wire_82, {c3540_wire_82_0, c3540_wire_82_1, c3540_wire_82_2, c3540_wire_82_3, c3540_wire_82_4});
fanout_n #(6, 0, 0) FANOUT_72 (c3540_wire_83, {c3540_wire_83_0, c3540_wire_83_1, c3540_wire_83_2, c3540_wire_83_3, c3540_wire_83_4, c3540_wire_83_5});
fanout_n #(4, 0, 0) FANOUT_73 (c3540_wire_84, {c3540_wire_84_0, c3540_wire_84_1, c3540_wire_84_2, c3540_wire_84_3});
fanout_n #(4, 0, 0) FANOUT_74 (c3540_wire_782, {c3540_wire_782_0, c3540_wire_782_1, c3540_wire_782_2, c3540_wire_782_3});
fanout_n #(2, 0, 0) FANOUT_75 (c3540_wire_159, {c3540_wire_159_0, c3540_wire_159_1});
fanout_n #(13, 0, 0) FANOUT_76 (c3540_wire_149, {c3540_wire_149_0, c3540_wire_149_1, c3540_wire_149_2, c3540_wire_149_3, c3540_wire_149_4, c3540_wire_149_5, c3540_wire_149_6, c3540_wire_149_7, c3540_wire_149_8, c3540_wire_149_9, c3540_wire_149_10, c3540_wire_149_11, c3540_wire_149_12});
fanout_n #(3, 0, 0) FANOUT_77 (c3540_wire_740, {c3540_wire_740_0, c3540_wire_740_1, c3540_wire_740_2});
fanout_n #(6, 0, 0) FANOUT_78 (c3540_wire_85, {c3540_wire_85_0, c3540_wire_85_1, c3540_wire_85_2, c3540_wire_85_3, c3540_wire_85_4, c3540_wire_85_5});
fanout_n #(2, 0, 0) FANOUT_79 (c3540_wire_158, {c3540_wire_158_0, c3540_wire_158_1});
fanout_n #(14, 0, 0) FANOUT_80 (c3540_wire_151, {c3540_wire_151_0, c3540_wire_151_1, c3540_wire_151_2, c3540_wire_151_3, c3540_wire_151_4, c3540_wire_151_5, c3540_wire_151_6, c3540_wire_151_7, c3540_wire_151_8, c3540_wire_151_9, c3540_wire_151_10, c3540_wire_151_11, c3540_wire_151_12, c3540_wire_151_13});
fanout_n #(2, 0, 0) FANOUT_81 (c3540_wire_805, {c3540_wire_805_0, c3540_wire_805_1});
fanout_n #(3, 0, 0) FANOUT_82 (c3540_wire_807, {c3540_wire_807_0, c3540_wire_807_1, c3540_wire_807_2});
fanout_n #(10, 0, 0) FANOUT_83 (c3540_wire_815, {c3540_wire_815_0, c3540_wire_815_1, c3540_wire_815_2, c3540_wire_815_3, c3540_wire_815_4, c3540_wire_815_5, c3540_wire_815_6, c3540_wire_815_7, c3540_wire_815_8, c3540_wire_815_9});
fanout_n #(7, 0, 0) FANOUT_84 (c3540_wire_827, {c3540_wire_827_0, c3540_wire_827_1, c3540_wire_827_2, c3540_wire_827_3, c3540_wire_827_4, c3540_wire_827_5, c3540_wire_827_6});
fanout_n #(6, 0, 0) FANOUT_85 (c3540_wire_41, {c3540_wire_41_0, c3540_wire_41_1, c3540_wire_41_2, c3540_wire_41_3, c3540_wire_41_4, c3540_wire_41_5});
fanout_n #(2, 0, 0) FANOUT_86 (c3540_wire_836, {c3540_wire_836_0, c3540_wire_836_1});
fanout_n #(10, 0, 0) FANOUT_87 (c3540_wire_799, {c3540_wire_799_0, c3540_wire_799_1, c3540_wire_799_2, c3540_wire_799_3, c3540_wire_799_4, c3540_wire_799_5, c3540_wire_799_6, c3540_wire_799_7, c3540_wire_799_8, c3540_wire_799_9});
fanout_n #(9, 0, 0) FANOUT_88 (c3540_wire_800, {c3540_wire_800_0, c3540_wire_800_1, c3540_wire_800_2, c3540_wire_800_3, c3540_wire_800_4, c3540_wire_800_5, c3540_wire_800_6, c3540_wire_800_7, c3540_wire_800_8});
fanout_n #(3, 0, 0) FANOUT_89 (c3540_wire_855, {c3540_wire_855_0, c3540_wire_855_1, c3540_wire_855_2});
fanout_n #(7, 0, 0) FANOUT_90 (c3540_wire_785, {c3540_wire_785_0, c3540_wire_785_1, c3540_wire_785_2, c3540_wire_785_3, c3540_wire_785_4, c3540_wire_785_5, c3540_wire_785_6});
fanout_n #(8, 0, 0) FANOUT_91 (c3540_wire_864, {c3540_wire_864_0, c3540_wire_864_1, c3540_wire_864_2, c3540_wire_864_3, c3540_wire_864_4, c3540_wire_864_5, c3540_wire_864_6, c3540_wire_864_7});
fanout_n #(5, 0, 0) FANOUT_92 (c3540_wire_904, {c3540_wire_904_0, c3540_wire_904_1, c3540_wire_904_2, c3540_wire_904_3, c3540_wire_904_4});
fanout_n #(5, 0, 0) FANOUT_93 (c3540_wire_909, {c3540_wire_909_0, c3540_wire_909_1, c3540_wire_909_2, c3540_wire_909_3, c3540_wire_909_4});
fanout_n #(2, 0, 0) FANOUT_94 (c3540_wire_916, {c3540_wire_916_0, c3540_wire_916_1});
fanout_n #(2, 0, 0) FANOUT_95 (c3540_wire_917, {c3540_wire_917_0, c3540_wire_917_1});
fanout_n #(4, 0, 0) FANOUT_96 (c3540_wire_935, {c3540_wire_935_0, c3540_wire_935_1, c3540_wire_935_2, c3540_wire_935_3});
fanout_n #(2, 0, 0) FANOUT_97 (c3540_wire_938, {c3540_wire_938_0, c3540_wire_938_1});
fanout_n #(4, 0, 0) FANOUT_98 (c3540_wire_942, {c3540_wire_942_0, c3540_wire_942_1, c3540_wire_942_2, c3540_wire_942_3});
fanout_n #(2, 0, 0) FANOUT_99 (c3540_wire_940, {c3540_wire_940_0, c3540_wire_940_1});
fanout_n #(2, 0, 0) FANOUT_100 (c3540_wire_333, {c3540_wire_333_0, c3540_wire_333_1});
fanout_n #(4, 0, 0) FANOUT_101 (c3540_wire_943, {c3540_wire_943_0, c3540_wire_943_1, c3540_wire_943_2, c3540_wire_943_3});
fanout_n #(3, 0, 0) FANOUT_102 (c3540_wire_946, {c3540_wire_946_0, c3540_wire_946_1, c3540_wire_946_2});
fanout_n #(2, 0, 0) FANOUT_103 (c3540_wire_952, {c3540_wire_952_0, c3540_wire_952_1});
fanout_n #(4, 0, 0) FANOUT_104 (c3540_wire_913, {c3540_wire_913_0, c3540_wire_913_1, c3540_wire_913_2, c3540_wire_913_3});
fanout_n #(2, 0, 0) FANOUT_105 (c3540_wire_837, {c3540_wire_837_0, c3540_wire_837_1});
fanout_n #(2, 0, 0) FANOUT_106 (c3540_wire_958, {c3540_wire_958_0, c3540_wire_958_1});
fanout_n #(40, 0, 0) FANOUT_107 (c3540_wire_33, {c3540_wire_33_0, c3540_wire_33_1, c3540_wire_33_2, c3540_wire_33_3, c3540_wire_33_4, c3540_wire_33_5, c3540_wire_33_6, c3540_wire_33_7, c3540_wire_33_8, c3540_wire_33_9, c3540_wire_33_10, c3540_wire_33_11, c3540_wire_33_12, c3540_wire_33_13, c3540_wire_33_14, c3540_wire_33_15, c3540_wire_33_16, c3540_wire_33_17, c3540_wire_33_18, c3540_wire_33_19, c3540_wire_33_20, c3540_wire_33_21, c3540_wire_33_22, c3540_wire_33_23, c3540_wire_33_24, c3540_wire_33_25, c3540_wire_33_26, c3540_wire_33_27, c3540_wire_33_28, c3540_wire_33_29, c3540_wire_33_30, c3540_wire_33_31, c3540_wire_33_32, c3540_wire_33_33, c3540_wire_33_34, c3540_wire_33_35, c3540_wire_33_36, c3540_wire_33_37, c3540_wire_33_38, c3540_wire_33_39});
fanout_n #(6, 0, 0) FANOUT_108 (c3540_wire_9, {c3540_wire_9_0, c3540_wire_9_1, c3540_wire_9_2, c3540_wire_9_3, c3540_wire_9_4, c3540_wire_9_5});
fanout_n #(4, 0, 0) FANOUT_109 (c3540_wire_973, {c3540_wire_973_0, c3540_wire_973_1, c3540_wire_973_2, c3540_wire_973_3});
fanout_n #(6, 0, 0) FANOUT_110 (c3540_wire_10, {c3540_wire_10_0, c3540_wire_10_1, c3540_wire_10_2, c3540_wire_10_3, c3540_wire_10_4, c3540_wire_10_5});
fanout_n #(5, 0, 0) FANOUT_111 (c3540_wire_1019, {c3540_wire_1019_0, c3540_wire_1019_1, c3540_wire_1019_2, c3540_wire_1019_3, c3540_wire_1019_4});
fanout_n #(4, 0, 0) FANOUT_112 (c3540_wire_1023, {c3540_wire_1023_0, c3540_wire_1023_1, c3540_wire_1023_2, c3540_wire_1023_3});
fanout_n #(4, 0, 0) FANOUT_113 (c3540_wire_1028, {c3540_wire_1028_0, c3540_wire_1028_1, c3540_wire_1028_2, c3540_wire_1028_3});
fanout_n #(2, 0, 0) FANOUT_114 (c3540_wire_1030, {c3540_wire_1030_0, c3540_wire_1030_1});
fanout_n #(5, 0, 0) FANOUT_115 (c3540_wire_824, {c3540_wire_824_0, c3540_wire_824_1, c3540_wire_824_2, c3540_wire_824_3, c3540_wire_824_4});
fanout_n #(4, 0, 0) FANOUT_116 (c3540_wire_1045, {c3540_wire_1045_0, c3540_wire_1045_1, c3540_wire_1045_2, c3540_wire_1045_3});
fanout_n #(8, 0, 0) FANOUT_117 (c3540_wire_401, {c3540_wire_401_0, c3540_wire_401_1, c3540_wire_401_2, c3540_wire_401_3, c3540_wire_401_4, c3540_wire_401_5, c3540_wire_401_6, c3540_wire_401_7});
fanout_n #(5, 0, 0) FANOUT_118 (c3540_wire_976, {c3540_wire_976_0, c3540_wire_976_1, c3540_wire_976_2, c3540_wire_976_3, c3540_wire_976_4});
fanout_n #(7, 0, 0) FANOUT_119 (c3540_wire_1104, {c3540_wire_1104_0, c3540_wire_1104_1, c3540_wire_1104_2, c3540_wire_1104_3, c3540_wire_1104_4, c3540_wire_1104_5, c3540_wire_1104_6});
fanout_n #(5, 0, 0) FANOUT_120 (c3540_wire_1122, {c3540_wire_1122_0, c3540_wire_1122_1, c3540_wire_1122_2, c3540_wire_1122_3, c3540_wire_1122_4});
fanout_n #(7, 0, 0) FANOUT_121 (c3540_wire_1159, {c3540_wire_1159_0, c3540_wire_1159_1, c3540_wire_1159_2, c3540_wire_1159_3, c3540_wire_1159_4, c3540_wire_1159_5, c3540_wire_1159_6});
fanout_n #(8, 0, 0) FANOUT_122 (c3540_wire_430, {c3540_wire_430_0, c3540_wire_430_1, c3540_wire_430_2, c3540_wire_430_3, c3540_wire_430_4, c3540_wire_430_5, c3540_wire_430_6, c3540_wire_430_7});
fanout_n #(6, 0, 0) FANOUT_123 (c3540_wire_1167, {c3540_wire_1167_0, c3540_wire_1167_1, c3540_wire_1167_2, c3540_wire_1167_3, c3540_wire_1167_4, c3540_wire_1167_5});
fanout_n #(4, 0, 0) FANOUT_124 (c3540_wire_1173, {c3540_wire_1173_0, c3540_wire_1173_1, c3540_wire_1173_2, c3540_wire_1173_3});
fanout_n #(6, 0, 0) FANOUT_125 (c3540_wire_1180, {c3540_wire_1180_0, c3540_wire_1180_1, c3540_wire_1180_2, c3540_wire_1180_3, c3540_wire_1180_4, c3540_wire_1180_5});
fanout_n #(2, 0, 0) FANOUT_126 (c3540_wire_1186, {c3540_wire_1186_0, c3540_wire_1186_1});
fanout_n #(7, 0, 0) FANOUT_127 (c3540_wire_28, {c3540_wire_28_0, c3540_wire_28_1, c3540_wire_28_2, c3540_wire_28_3, c3540_wire_28_4, c3540_wire_28_5, c3540_wire_28_6});
fanout_n #(2, 0, 0) FANOUT_128 (c3540_wire_1193, {c3540_wire_1193_0, c3540_wire_1193_1});
fanout_n #(4, 0, 0) FANOUT_129 (c3540_wire_1195, {c3540_wire_1195_0, c3540_wire_1195_1, c3540_wire_1195_2, c3540_wire_1195_3});
fanout_n #(2, 0, 0) FANOUT_130 (c3540_wire_1196, {c3540_wire_1196_0, c3540_wire_1196_1});
fanout_n #(3, 0, 0) FANOUT_131 (c3540_wire_1200, {c3540_wire_1200_0, c3540_wire_1200_1, c3540_wire_1200_2});
fanout_n #(7, 0, 0) FANOUT_132 (c3540_wire_111, {c3540_wire_111_0, c3540_wire_111_1, c3540_wire_111_2, c3540_wire_111_3, c3540_wire_111_4, c3540_wire_111_5, c3540_wire_111_6});
fanout_n #(6, 0, 0) FANOUT_133 (c3540_wire_115, {c3540_wire_115_0, c3540_wire_115_1, c3540_wire_115_2, c3540_wire_115_3, c3540_wire_115_4, c3540_wire_115_5});
fanout_n #(4, 0, 0) FANOUT_134 (c3540_wire_116, {c3540_wire_116_0, c3540_wire_116_1, c3540_wire_116_2, c3540_wire_116_3});
fanout_n #(8, 0, 0) FANOUT_135 (c3540_wire_340, {c3540_wire_340_0, c3540_wire_340_1, c3540_wire_340_2, c3540_wire_340_3, c3540_wire_340_4, c3540_wire_340_5, c3540_wire_340_6, c3540_wire_340_7});
fanout_n #(9, 0, 0) FANOUT_136 (c3540_wire_483, {c3540_wire_483_0, c3540_wire_483_1, c3540_wire_483_2, c3540_wire_483_3, c3540_wire_483_4, c3540_wire_483_5, c3540_wire_483_6, c3540_wire_483_7, c3540_wire_483_8});
fanout_n #(4, 0, 0) FANOUT_137 (c3540_wire_326, {c3540_wire_326_0, c3540_wire_326_1, c3540_wire_326_2, c3540_wire_326_3});
fanout_n #(55, 0, 0) FANOUT_138 (c3540_wire_60, {c3540_wire_60_0, c3540_wire_60_1, c3540_wire_60_2, c3540_wire_60_3, c3540_wire_60_4, c3540_wire_60_5, c3540_wire_60_6, c3540_wire_60_7, c3540_wire_60_8, c3540_wire_60_9, c3540_wire_60_10, c3540_wire_60_11, c3540_wire_60_12, c3540_wire_60_13, c3540_wire_60_14, c3540_wire_60_15, c3540_wire_60_16, c3540_wire_60_17, c3540_wire_60_18, c3540_wire_60_19, c3540_wire_60_20, c3540_wire_60_21, c3540_wire_60_22, c3540_wire_60_23, c3540_wire_60_24, c3540_wire_60_25, c3540_wire_60_26, c3540_wire_60_27, c3540_wire_60_28, c3540_wire_60_29, c3540_wire_60_30, c3540_wire_60_31, c3540_wire_60_32, c3540_wire_60_33, c3540_wire_60_34, c3540_wire_60_35, c3540_wire_60_36, c3540_wire_60_37, c3540_wire_60_38, c3540_wire_60_39, c3540_wire_60_40, c3540_wire_60_41, c3540_wire_60_42, c3540_wire_60_43, c3540_wire_60_44, c3540_wire_60_45, c3540_wire_60_46, c3540_wire_60_47, c3540_wire_60_48, c3540_wire_60_49, c3540_wire_60_50, c3540_wire_60_51, c3540_wire_60_52, c3540_wire_60_53, c3540_wire_60_54});
fanout_n #(7, 0, 0) FANOUT_139 (c3540_wire_516, {c3540_wire_516_0, c3540_wire_516_1, c3540_wire_516_2, c3540_wire_516_3, c3540_wire_516_4, c3540_wire_516_5, c3540_wire_516_6});
fanout_n #(7, 0, 0) FANOUT_140 (c3540_wire_549, {c3540_wire_549_0, c3540_wire_549_1, c3540_wire_549_2, c3540_wire_549_3, c3540_wire_549_4, c3540_wire_549_5, c3540_wire_549_6});
fanout_n #(5, 0, 0) FANOUT_141 (c3540_wire_685, {c3540_wire_685_0, c3540_wire_685_1, c3540_wire_685_2, c3540_wire_685_3, c3540_wire_685_4});
fanout_n #(4, 0, 0) FANOUT_142 (c3540_wire_1002, {c3540_wire_1002_0, c3540_wire_1002_1, c3540_wire_1002_2, c3540_wire_1002_3});
fanout_n #(3, 0, 0) FANOUT_143 (c3540_wire_994, {c3540_wire_994_0, c3540_wire_994_1, c3540_wire_994_2});
fanout_n #(2, 0, 0) FANOUT_144 (c3540_wire_997, {c3540_wire_997_0, c3540_wire_997_1});
fanout_n #(15, 0, 0) FANOUT_145 (c3540_wire_832, {c3540_wire_832_0, c3540_wire_832_1, c3540_wire_832_2, c3540_wire_832_3, c3540_wire_832_4, c3540_wire_832_5, c3540_wire_832_6, c3540_wire_832_7, c3540_wire_832_8, c3540_wire_832_9, c3540_wire_832_10, c3540_wire_832_11, c3540_wire_832_12, c3540_wire_832_13, c3540_wire_832_14});
fanout_n #(2, 0, 0) FANOUT_146 (c3540_wire_42, {c3540_wire_42_0, c3540_wire_42_1});
fanout_n #(8, 0, 0) FANOUT_147 (c3540_wire_344, {c3540_wire_344_0, c3540_wire_344_1, c3540_wire_344_2, c3540_wire_344_3, c3540_wire_344_4, c3540_wire_344_5, c3540_wire_344_6, c3540_wire_344_7});
fanout_n #(4, 0, 0) FANOUT_148 (c3540_wire_449, {c3540_wire_449_0, c3540_wire_449_1, c3540_wire_449_2, c3540_wire_449_3});
fanout_n #(17, 0, 0) FANOUT_149 (c3540_wire_38, {c3540_wire_38_0, c3540_wire_38_1, c3540_wire_38_2, c3540_wire_38_3, c3540_wire_38_4, c3540_wire_38_5, c3540_wire_38_6, c3540_wire_38_7, c3540_wire_38_8, c3540_wire_38_9, c3540_wire_38_10, c3540_wire_38_11, c3540_wire_38_12, c3540_wire_38_13, c3540_wire_38_14, c3540_wire_38_15, c3540_wire_38_16});
fanout_n #(12, 0, 0) FANOUT_150 (c3540_wire_469, {c3540_wire_469_0, c3540_wire_469_1, c3540_wire_469_2, c3540_wire_469_3, c3540_wire_469_4, c3540_wire_469_5, c3540_wire_469_6, c3540_wire_469_7, c3540_wire_469_8, c3540_wire_469_9, c3540_wire_469_10, c3540_wire_469_11});
fanout_n #(5, 0, 0) FANOUT_151 (c3540_wire_1049, {c3540_wire_1049_0, c3540_wire_1049_1, c3540_wire_1049_2, c3540_wire_1049_3, c3540_wire_1049_4});
fanout_n #(19, 0, 0) FANOUT_152 (c3540_wire_18, {c3540_wire_18_0, c3540_wire_18_1, c3540_wire_18_2, c3540_wire_18_3, c3540_wire_18_4, c3540_wire_18_5, c3540_wire_18_6, c3540_wire_18_7, c3540_wire_18_8, c3540_wire_18_9, c3540_wire_18_10, c3540_wire_18_11, c3540_wire_18_12, c3540_wire_18_13, c3540_wire_18_14, c3540_wire_18_15, c3540_wire_18_16, c3540_wire_18_17, c3540_wire_18_18});
fanout_n #(2, 0, 0) FANOUT_153 (c3540_wire_309, {c3540_wire_309_0, c3540_wire_309_1});
fanout_n #(8, 0, 0) FANOUT_154 (c3540_wire_341, {c3540_wire_341_0, c3540_wire_341_1, c3540_wire_341_2, c3540_wire_341_3, c3540_wire_341_4, c3540_wire_341_5, c3540_wire_341_6, c3540_wire_341_7});
fanout_n #(3, 0, 0) FANOUT_155 (c3540_wire_492, {c3540_wire_492_0, c3540_wire_492_1, c3540_wire_492_2});
fanout_n #(19, 0, 0) FANOUT_156 (c3540_wire_120, {c3540_wire_120_0, c3540_wire_120_1, c3540_wire_120_2, c3540_wire_120_3, c3540_wire_120_4, c3540_wire_120_5, c3540_wire_120_6, c3540_wire_120_7, c3540_wire_120_8, c3540_wire_120_9, c3540_wire_120_10, c3540_wire_120_11, c3540_wire_120_12, c3540_wire_120_13, c3540_wire_120_14, c3540_wire_120_15, c3540_wire_120_16, c3540_wire_120_17, c3540_wire_120_18});
fanout_n #(16, 0, 0) FANOUT_157 (c3540_wire_318, {c3540_wire_318_0, c3540_wire_318_1, c3540_wire_318_2, c3540_wire_318_3, c3540_wire_318_4, c3540_wire_318_5, c3540_wire_318_6, c3540_wire_318_7, c3540_wire_318_8, c3540_wire_318_9, c3540_wire_318_10, c3540_wire_318_11, c3540_wire_318_12, c3540_wire_318_13, c3540_wire_318_14, c3540_wire_318_15});
fanout_n #(23, 0, 0) FANOUT_158 (c3540_wire_121, {c3540_wire_121_0, c3540_wire_121_1, c3540_wire_121_2, c3540_wire_121_3, c3540_wire_121_4, c3540_wire_121_5, c3540_wire_121_6, c3540_wire_121_7, c3540_wire_121_8, c3540_wire_121_9, c3540_wire_121_10, c3540_wire_121_11, c3540_wire_121_12, c3540_wire_121_13, c3540_wire_121_14, c3540_wire_121_15, c3540_wire_121_16, c3540_wire_121_17, c3540_wire_121_18, c3540_wire_121_19, c3540_wire_121_20, c3540_wire_121_21, c3540_wire_121_22});
fanout_n #(8, 0, 0) FANOUT_159 (c3540_wire_1009, {c3540_wire_1009_0, c3540_wire_1009_1, c3540_wire_1009_2, c3540_wire_1009_3, c3540_wire_1009_4, c3540_wire_1009_5, c3540_wire_1009_6, c3540_wire_1009_7});
fanout_n #(8, 0, 0) FANOUT_160 (c3540_wire_346, {c3540_wire_346_0, c3540_wire_346_1, c3540_wire_346_2, c3540_wire_346_3, c3540_wire_346_4, c3540_wire_346_5, c3540_wire_346_6, c3540_wire_346_7});


bufg #(0, 0) BUF_1 (c3540_wire_1, G1_net_0);
bufg #(0, 0) BUF_2 (c3540_wire_2, G10_net_0);
and_n #(2, 0, 0) AND_1 (c3540_wire_3, {c3540_wire_4, c3540_wire_5_0});
notg #(0, 0) NOT_1 (c3540_wire_6, c3540_wire_3);
notg #(0, 0) NOT_2 (c3540_wire_4, c3540_wire_7);
and_n #(2, 0, 0) AND_2 (c3540_wire_8, {c3540_wire_9_0, c3540_wire_10_0});
or_n #(2, 0, 0) OR_1 (c3540_wire_11, {c3540_wire_8, c3540_wire_12});
nor_n #(2, 0, 0) NOR_1 (c3540_wire_12, {c3540_wire_10_1, c3540_wire_9_1});
and_n #(2, 0, 0) AND_3 (c3540_wire_13, {c3540_wire_14, c3540_wire_15});
notg #(0, 0) NOT_3 (c3540_wire_16, c3540_wire_9_2);
or_n #(2, 0, 0) OR_2 (c3540_wire_17, {c3540_wire_16, c3540_wire_18_0});
or_n #(2, 0, 0) OR_3 (c3540_wire_19, {c3540_wire_20, c3540_wire_5_1});
and_n #(3, 0, 0) AND_4 (c3540_wire_15, {c3540_wire_19, c3540_wire_21, c3540_wire_17});
nor_n #(2, 0, 0) NOR_2 (c3540_wire_21, {c3540_wire_22, c3540_wire_23});
nor_n #(4, 0, 0) NOR_3 (c3540_wire_14, {c3540_wire_24, c3540_wire_25, c3540_wire_26, c3540_wire_27});
notg #(0, 0) NOT_4 (c3540_wire_20, c3540_wire_28_0);
notg #(0, 0) NOT_5 (c3540_wire_29, c3540_wire_1_0);
and_n #(3, 0, 0) AND_5 (c3540_wire_30, {c3540_wire_29, c3540_wire_31, c3540_wire_32_0});
notg #(0, 0) NOT_6 (c3540_wire_31, c3540_wire_33_0);
notg #(0, 0) NOT_7 (c3540_wire_34, c3540_wire_1_1);
and_n #(4, 0, 0) AND_6 (c3540_wire_35, {c3540_wire_34, c3540_wire_36, c3540_wire_37, c3540_wire_38_0});
notg #(0, 0) NOT_8 (c3540_wire_36, c3540_wire_32_1);
notg #(0, 0) NOT_9 (c3540_wire_37, c3540_wire_33_1);
nor_n #(3, 0, 0) NOR_4 (c3540_wire_39, {c3540_wire_32_2, c3540_wire_1_2, c3540_wire_33_2});
and_n #(3, 0, 0) AND_7 (c3540_wire_40, {c3540_wire_39_0, c3540_wire_41_0, c3540_wire_42_0});
and_n #(2, 0, 0) AND_8 (c3540_wire_43, {c3540_wire_39_1, c3540_wire_28_1});
and_n #(3, 0, 0) AND_9 (c3540_wire_44, {c3540_wire_39_2, c3540_wire_45_0, c3540_wire_41_1});
and_n #(3, 0, 0) AND_10 (c3540_wire_46, {c3540_wire_39_3, c3540_wire_47_0, c3540_wire_41_2});
and_n #(2, 0, 0) AND_11 (c3540_wire_48, {c3540_wire_39_4, c3540_wire_41_3});
notg #(0, 0) NOT_10 (c3540_wire_49, c3540_wire_2_0);
notg #(0, 0) NOT_11 (c3540_wire_50, c3540_wire_2_1);
notg #(0, 0) NOT_12 (c3540_wire_51, c3540_wire_2_2);
and_n #(2, 0, 0) AND_12 (c3540_wire_52, {c3540_wire_2_3, c3540_wire_53});
or_n #(2, 0, 0) OR_4 (c3540_wire_54, {c3540_wire_2_4, c3540_wire_55});
notg #(0, 0) NOT_13 (c3540_wire_56, c3540_wire_2_5);
and_n #(2, 0, 0) AND_13 (c3540_wire_57, {c3540_wire_2_6, c3540_wire_58});
and_n #(2, 0, 0) AND_14 (c3540_wire_59, {c3540_wire_2_7, c3540_wire_60_0});
and_n #(2, 0, 0) AND_15 (c3540_wire_61, {c3540_wire_2_8, c3540_wire_62});
notg #(0, 0) NOT_14 (c3540_wire_63, c3540_wire_2_9);
notg #(0, 0) NOT_15 (c3540_wire_64, c3540_wire_2_10);
notg #(0, 0) NOT_16 (c3540_wire_65, c3540_wire_2_11);
bufg #(0, 0) BUF_3 (c3540_wire_5, G11_net_0);
notg #(0, 0) NOT_17 (c3540_wire_66, c3540_wire_40_0);
notg #(0, 0) NOT_18 (c3540_wire_67, c3540_wire_40_1);
and_n #(2, 0, 0) AND_16 (c3540_wire_68, {c3540_wire_40_2, c3540_wire_69_0});
and_n #(2, 0, 0) AND_17 (c3540_wire_70, {c3540_wire_40_3, c3540_wire_71_0});
and_n #(2, 0, 0) AND_18 (c3540_wire_72, {c3540_wire_40_4, c3540_wire_73_0});
and_n #(2, 0, 0) AND_19 (c3540_wire_74, {c3540_wire_40_5, c3540_wire_75_0});
and_n #(2, 0, 0) AND_20 (c3540_wire_76, {c3540_wire_40_6, c3540_wire_77_0});
and_n #(2, 0, 0) AND_21 (c3540_wire_78, {c3540_wire_40_7, c3540_wire_79_0});
notg #(0, 0) NOT_19 (c3540_wire_80, c3540_wire_40_8);
and_n #(5, 0, 0) AND_22 (c3540_wire_81, {c3540_wire_40_9, c3540_wire_82_0, c3540_wire_83_0, c3540_wire_84_0, c3540_wire_85_0});
notg #(0, 0) NOT_20 (c3540_wire_86, c3540_wire_40_10);
or_n #(2, 0, 0) OR_5 (c3540_wire_87, {c3540_wire_40_11, c3540_wire_88});
notg #(0, 0) NOT_21 (c3540_wire_89, c3540_wire_40_12);
notg #(0, 0) NOT_22 (c3540_wire_90, c3540_wire_40_13);
or_n #(2, 0, 0) OR_6 (c3540_wire_91, {c3540_wire_40_14, c3540_wire_92});
and_n #(2, 0, 0) AND_23 (c3540_wire_93, {c3540_wire_41_4, c3540_wire_42_1});
notg #(0, 0) NOT_23 (c3540_wire_94, c3540_wire_93_0);
notg #(0, 0) NOT_24 (c3540_wire_95, c3540_wire_93_1);
or_n #(2, 0, 0) OR_7 (c3540_wire_96, {c3540_wire_93_2, c3540_wire_97});
and_n #(2, 0, 0) AND_24 (c3540_wire_98, {c3540_wire_5_2, c3540_wire_99_0});
notg #(0, 0) NOT_25 (c3540_wire_100, c3540_wire_5_3);
notg #(0, 0) NOT_26 (c3540_wire_101, c3540_wire_5_4);
or_n #(2, 0, 0) OR_8 (c3540_wire_102, {c3540_wire_5_5, c3540_wire_103});
notg #(0, 0) NOT_27 (c3540_wire_104, c3540_wire_5_6);
notg #(0, 0) NOT_28 (c3540_wire_105, c3540_wire_5_7);
and_n #(4, 0, 0) AND_25 (c3540_wire_106, {c3540_wire_5_8, c3540_wire_107, c3540_wire_108, c3540_wire_109});
bufg #(0, 0) BUF_4 (c3540_wire_99, G12_net_0);
and_n #(2, 0, 0) AND_26 (c3540_wire_110, {c3540_wire_28_2, c3540_wire_111_0});
or_n #(2, 0, 0) OR_9 (c3540_wire_112, {c3540_wire_110, c3540_wire_113});
nor_n #(2, 0, 0) NOR_5 (c3540_wire_113, {c3540_wire_111_1, c3540_wire_28_3});
and_n #(2, 0, 0) AND_27 (c3540_wire_114, {c3540_wire_115_0, c3540_wire_116_0});
or_n #(2, 0, 0) OR_10 (c3540_wire_117, {c3540_wire_114, c3540_wire_118});
nor_n #(2, 0, 0) NOR_6 (c3540_wire_118, {c3540_wire_116_1, c3540_wire_115_1});
nor_n #(2, 0, 0) NOR_7 (c3540_wire_119, {c3540_wire_120_0, c3540_wire_121_0});
notg #(0, 0) NOT_29 (c3540_wire_122, c3540_wire_119_0);
nor_n #(2, 0, 0) NOR_8 (c3540_wire_7, {c3540_wire_99_1, c3540_wire_123_0});
notg #(0, 0) NOT_30 (c3540_wire_124, c3540_wire_99_2);
xor_n #(2, 0, 0) XOR_1 (c3540_wire_125, {c3540_wire_99_3, c3540_wire_123_1});
notg #(0, 0) NOT_31 (c3540_wire_126, c3540_wire_99_4);
or_n #(2, 0, 0) OR_11 (c3540_wire_127, {c3540_wire_99_5, c3540_wire_128});
notg #(0, 0) NOT_32 (c3540_wire_129, c3540_wire_99_6);
notg #(0, 0) NOT_33 (c3540_wire_130, c3540_wire_99_7);
and_n #(4, 0, 0) AND_28 (c3540_wire_131, {c3540_wire_99_8, c3540_wire_132, c3540_wire_133, c3540_wire_134});
notg #(0, 0) NOT_34 (c3540_wire_135, c3540_wire_99_9);
bufg #(0, 0) BUF_5 (c3540_wire_123, G13_net_0);
and_n #(2, 0, 0) AND_29 (c3540_wire_136, {c3540_wire_112_0, c3540_wire_137});
xor_n #(2, 0, 0) XOR_2 (c3540_wire_137, {c3540_wire_117_0, c3540_wire_138_0});
xor_n #(2, 0, 0) XOR_3 (c3540_wire_139, {c3540_wire_117_1, c3540_wire_138_1});
notg #(0, 0) NOT_35 (c3540_wire_140, c3540_wire_35_0);
notg #(0, 0) NOT_36 (c3540_wire_141, c3540_wire_35_1);
notg #(0, 0) NOT_37 (c3540_wire_142, c3540_wire_35_2);
notg #(0, 0) NOT_38 (c3540_wire_143, c3540_wire_35_3);
notg #(0, 0) NOT_39 (c3540_wire_144, c3540_wire_35_4);
notg #(0, 0) NOT_40 (c3540_wire_145, c3540_wire_35_5);
and_n #(3, 0, 0) AND_30 (c3540_wire_146, {c3540_wire_30_0, c3540_wire_122, c3540_wire_147});
nor_n #(3, 0, 0) NOR_9 (c3540_wire_148, {c3540_wire_149_0, c3540_wire_150_0, c3540_wire_151_0});
notg #(0, 0) NOT_41 (c3540_wire_152, c3540_wire_33_3);
or_n #(2, 0, 0) OR_12 (c3540_wire_153, {c3540_wire_152, c3540_wire_148});
and_n #(2, 0, 0) AND_31 (c3540_wire_154, {c3540_wire_151_1, c3540_wire_33_4});
and_n #(2, 0, 0) AND_32 (c3540_wire_155, {c3540_wire_154, c3540_wire_156});
nor_n #(2, 0, 0) NOR_10 (c3540_wire_156, {c3540_wire_149_1, c3540_wire_150_1});
nor_n #(3, 0, 0) NOR_11 (c3540_wire_157, {c3540_wire_151_2, c3540_wire_158_0, c3540_wire_159_0});
notg #(0, 0) NOT_42 (c3540_wire_160, c3540_wire_158_1);
and_n #(3, 0, 0) AND_33 (c3540_wire_161, {c3540_wire_160, c3540_wire_162, c3540_wire_151_3});
notg #(0, 0) NOT_43 (c3540_wire_162, c3540_wire_159_1);
and_n #(3, 0, 0) AND_34 (c3540_wire_163, {c3540_wire_164, c3540_wire_165, c3540_wire_32_3});
notg #(0, 0) NOT_44 (c3540_wire_166, c3540_wire_163_0);
and_n #(2, 0, 0) AND_35 (c3540_wire_167, {c3540_wire_163_1, c3540_wire_168});
notg #(0, 0) NOT_45 (c3540_wire_169, c3540_wire_163_2);
and_n #(2, 0, 0) AND_36 (c3540_wire_170, {c3540_wire_163_3, c3540_wire_171});
notg #(0, 0) NOT_46 (c3540_wire_172, c3540_wire_163_4);
and_n #(2, 0, 0) AND_37 (c3540_wire_173, {c3540_wire_163_5, c3540_wire_51});
notg #(0, 0) NOT_47 (c3540_wire_174, c3540_wire_163_6);
and_n #(2, 0, 0) AND_38 (c3540_wire_175, {c3540_wire_163_7, c3540_wire_176});
notg #(0, 0) NOT_48 (c3540_wire_177, c3540_wire_33_5);
or_n #(2, 0, 0) OR_13 (c3540_wire_165, {c3540_wire_177, c3540_wire_178_0});
notg #(0, 0) NOT_49 (c3540_wire_164, c3540_wire_1_3);
notg #(0, 0) NOT_50 (c3540_wire_179, c3540_wire_123_2);
and_n #(2, 0, 0) AND_39 (c3540_wire_180, {c3540_wire_123_3, c3540_wire_181_0});
notg #(0, 0) NOT_51 (c3540_wire_182, c3540_wire_123_4);
or_n #(2, 0, 0) OR_14 (c3540_wire_183, {c3540_wire_123_5, c3540_wire_184});
notg #(0, 0) NOT_52 (c3540_wire_185, c3540_wire_123_6);
and_n #(4, 0, 0) AND_40 (c3540_wire_186, {c3540_wire_123_7, c3540_wire_187, c3540_wire_188, c3540_wire_189});
and_n #(2, 0, 0) AND_41 (c3540_wire_190, {c3540_wire_123_8, c3540_wire_60_1});
notg #(0, 0) NOT_53 (c3540_wire_191, c3540_wire_123_9);
bufg #(0, 0) BUF_6 (c3540_wire_181, G14_net_0);
and_n #(2, 0, 0) AND_42 (c3540_wire_192, {c3540_wire_94, c3540_wire_193});
and_n #(2, 0, 0) AND_43 (c3540_wire_194, {c3540_wire_192_0, c3540_wire_195});
and_n #(2, 0, 0) AND_44 (c3540_wire_196, {c3540_wire_11_0, c3540_wire_197});
or_n #(2, 0, 0) OR_15 (c3540_wire_198, {c3540_wire_98, c3540_wire_199});
nor_n #(2, 0, 0) NOR_12 (c3540_wire_199, {c3540_wire_99_10, c3540_wire_5_9});
or_n #(2, 0, 0) OR_16 (c3540_wire_200, {c3540_wire_180, c3540_wire_201});
nor_n #(2, 0, 0) NOR_13 (c3540_wire_201, {c3540_wire_181_1, c3540_wire_123_10});
and_n #(2, 0, 0) AND_45 (c3540_wire_202, {c3540_wire_125_0, c3540_wire_33_6});
notg #(0, 0) NOT_54 (c3540_wire_203, c3540_wire_125_1);
notg #(0, 0) NOT_55 (c3540_wire_204, c3540_wire_181_2);
notg #(0, 0) NOT_56 (c3540_wire_205, c3540_wire_181_3);
or_n #(2, 0, 0) OR_17 (c3540_wire_206, {c3540_wire_181_4, c3540_wire_207});
notg #(0, 0) NOT_57 (c3540_wire_208, c3540_wire_181_5);
and_n #(2, 0, 0) AND_46 (c3540_wire_209, {c3540_wire_181_6, c3540_wire_210});
and_n #(2, 0, 0) AND_47 (c3540_wire_211, {c3540_wire_181_7, c3540_wire_60_2});
notg #(0, 0) NOT_58 (c3540_wire_212, c3540_wire_181_8);
notg #(0, 0) NOT_59 (c3540_wire_213, c3540_wire_181_9);
bufg #(0, 0) BUF_7 (c3540_wire_214, G15_net_0);
xor_n #(2, 0, 0) XOR_4 (c3540_wire_215, {c3540_wire_18_1, c3540_wire_120_1});
and_n #(2, 0, 0) AND_48 (c3540_wire_216, {c3540_wire_215_0, c3540_wire_121_1});
and_n #(2, 0, 0) AND_49 (c3540_wire_217, {c3540_wire_215_1, c3540_wire_121_2});
and_n #(2, 0, 0) AND_50 (c3540_wire_218, {c3540_wire_198_0, c3540_wire_219});
and_n #(2, 0, 0) AND_51 (c3540_wire_220, {c3540_wire_200_0, c3540_wire_221_0});
and_n #(2, 0, 0) AND_52 (c3540_wire_222, {c3540_wire_200_1, c3540_wire_221_1});
notg #(0, 0) NOT_60 (c3540_wire_223, c3540_wire_224_0);
notg #(0, 0) NOT_61 (c3540_wire_225, c3540_wire_224_1);
notg #(0, 0) NOT_62 (c3540_wire_226, c3540_wire_224_2);
notg #(0, 0) NOT_63 (c3540_wire_227, c3540_wire_224_3);
notg #(0, 0) NOT_64 (c3540_wire_228, c3540_wire_224_4);
notg #(0, 0) NOT_65 (c3540_wire_229, c3540_wire_224_5);
notg #(0, 0) NOT_66 (c3540_wire_230, c3540_wire_224_6);
notg #(0, 0) NOT_67 (c3540_wire_231, c3540_wire_224_7);
and_n #(2, 0, 0) AND_53 (c3540_wire_224, {c3540_wire_232, c3540_wire_233});
notg #(0, 0) NOT_68 (c3540_wire_234, c3540_wire_224_8);
notg #(0, 0) NOT_69 (c3540_wire_235, c3540_wire_224_9);
notg #(0, 0) NOT_70 (c3540_wire_236, c3540_wire_224_10);
notg #(0, 0) NOT_71 (c3540_wire_237, c3540_wire_224_11);
notg #(0, 0) NOT_72 (c3540_wire_238, c3540_wire_224_12);
notg #(0, 0) NOT_73 (c3540_wire_239, c3540_wire_224_13);
notg #(0, 0) NOT_74 (c3540_wire_240, c3540_wire_224_14);
notg #(0, 0) NOT_75 (c3540_wire_241, c3540_wire_224_15);
and_n #(2, 0, 0) AND_54 (c3540_wire_232, {c3540_wire_149_2, c3540_wire_33_7});
nor_n #(2, 0, 0) NOR_14 (c3540_wire_233, {c3540_wire_151_4, c3540_wire_150_2});
and_n #(2, 0, 0) AND_55 (c3540_wire_242, {c3540_wire_243, c3540_wire_244});
notg #(0, 0) NOT_76 (c3540_wire_245, c3540_wire_242_0);
notg #(0, 0) NOT_77 (c3540_wire_246, c3540_wire_242_1);
notg #(0, 0) NOT_78 (c3540_wire_247, c3540_wire_242_2);
notg #(0, 0) NOT_79 (c3540_wire_248, c3540_wire_242_3);
notg #(0, 0) NOT_80 (c3540_wire_249, c3540_wire_242_4);
notg #(0, 0) NOT_81 (c3540_wire_250, c3540_wire_242_5);
notg #(0, 0) NOT_82 (c3540_wire_251, c3540_wire_242_6);
notg #(0, 0) NOT_83 (c3540_wire_252, c3540_wire_242_7);
notg #(0, 0) NOT_84 (c3540_wire_253, c3540_wire_242_8);
notg #(0, 0) NOT_85 (c3540_wire_254, c3540_wire_242_9);
notg #(0, 0) NOT_86 (c3540_wire_255, c3540_wire_242_10);
notg #(0, 0) NOT_87 (c3540_wire_256, c3540_wire_242_11);
notg #(0, 0) NOT_88 (c3540_wire_257, c3540_wire_242_12);
notg #(0, 0) NOT_89 (c3540_wire_258, c3540_wire_242_13);
notg #(0, 0) NOT_90 (c3540_wire_259, c3540_wire_242_14);
notg #(0, 0) NOT_91 (c3540_wire_260, c3540_wire_242_15);
and_n #(2, 0, 0) AND_56 (c3540_wire_243, {c3540_wire_149_3, c3540_wire_33_8});
notg #(0, 0) NOT_92 (c3540_wire_261, c3540_wire_150_3);
and_n #(2, 0, 0) AND_57 (c3540_wire_244, {c3540_wire_261, c3540_wire_151_5});
notg #(0, 0) NOT_93 (c3540_wire_262, c3540_wire_153_0);
notg #(0, 0) NOT_94 (c3540_wire_263, c3540_wire_153_1);
notg #(0, 0) NOT_95 (c3540_wire_264, c3540_wire_155_0);
notg #(0, 0) NOT_96 (c3540_wire_265, c3540_wire_155_1);
notg #(0, 0) NOT_97 (c3540_wire_266, c3540_wire_155_2);
notg #(0, 0) NOT_98 (c3540_wire_267, c3540_wire_155_3);
notg #(0, 0) NOT_99 (c3540_wire_268, c3540_wire_155_4);
notg #(0, 0) NOT_100 (c3540_wire_269, c3540_wire_155_5);
notg #(0, 0) NOT_101 (c3540_wire_270, c3540_wire_157_0);
notg #(0, 0) NOT_102 (c3540_wire_271, c3540_wire_157_1);
notg #(0, 0) NOT_103 (c3540_wire_272, c3540_wire_157_2);
notg #(0, 0) NOT_104 (c3540_wire_273, c3540_wire_157_3);
notg #(0, 0) NOT_105 (c3540_wire_274, c3540_wire_157_4);
notg #(0, 0) NOT_106 (c3540_wire_275, c3540_wire_157_5);
notg #(0, 0) NOT_107 (c3540_wire_276, c3540_wire_157_6);
notg #(0, 0) NOT_108 (c3540_wire_277, c3540_wire_157_7);
notg #(0, 0) NOT_109 (c3540_wire_278, c3540_wire_157_8);
notg #(0, 0) NOT_110 (c3540_wire_279, c3540_wire_157_9);
notg #(0, 0) NOT_111 (c3540_wire_280, c3540_wire_157_10);
notg #(0, 0) NOT_112 (c3540_wire_281, c3540_wire_157_11);
notg #(0, 0) NOT_113 (c3540_wire_282, c3540_wire_161_0);
notg #(0, 0) NOT_114 (c3540_wire_283, c3540_wire_161_1);
notg #(0, 0) NOT_115 (c3540_wire_284, c3540_wire_161_2);
notg #(0, 0) NOT_116 (c3540_wire_285, c3540_wire_161_3);
notg #(0, 0) NOT_117 (c3540_wire_286, c3540_wire_161_4);
notg #(0, 0) NOT_118 (c3540_wire_287, c3540_wire_161_5);
notg #(0, 0) NOT_119 (c3540_wire_288, c3540_wire_161_6);
notg #(0, 0) NOT_120 (c3540_wire_289, c3540_wire_161_7);
notg #(0, 0) NOT_121 (c3540_wire_290, c3540_wire_161_8);
notg #(0, 0) NOT_122 (c3540_wire_291, c3540_wire_161_9);
notg #(0, 0) NOT_123 (c3540_wire_292, c3540_wire_161_10);
notg #(0, 0) NOT_124 (c3540_wire_293, c3540_wire_161_11);
notg #(0, 0) NOT_125 (c3540_wire_294, c3540_wire_161_12);
notg #(0, 0) NOT_126 (c3540_wire_295, c3540_wire_161_13);
or_n #(2, 0, 0) OR_18 (c3540_wire_296, {c3540_wire_214, c3540_wire_297_0});
bufg #(0, 0) BUF_8 (c3540_wire_298, G16_net_0);
and_n #(3, 0, 0) AND_58 (c3540_wire_299, {c3540_wire_45_1, c3540_wire_300, c3540_wire_301});
notg #(0, 0) NOT_127 (c3540_wire_302, c3540_wire_45_2);
and_n #(2, 0, 0) AND_59 (c3540_wire_303, {c3540_wire_45_3, c3540_wire_304});
or_n #(3, 0, 0) OR_19 (c3540_wire_45, {c3540_wire_305, c3540_wire_306, c3540_wire_307});
notg #(0, 0) NOT_128 (c3540_wire_308, c3540_wire_309_0);
and_n #(2, 0, 0) AND_60 (c3540_wire_310, {c3540_wire_308, c3540_wire_33_9});
and_n #(2, 0, 0) AND_61 (c3540_wire_311, {c3540_wire_312, c3540_wire_313_0});
or_n #(2, 0, 0) OR_20 (c3540_wire_314, {c3540_wire_311, c3540_wire_315});
and_n #(2, 0, 0) AND_62 (c3540_wire_315, {c3540_wire_316, c3540_wire_60_3});
and_n #(2, 0, 0) AND_63 (c3540_wire_305, {c3540_wire_317, c3540_wire_318_0});
and_n #(4, 0, 0) AND_64 (c3540_wire_306, {c3540_wire_319, c3540_wire_320, c3540_wire_321, c3540_wire_18_2});
and_n #(2, 0, 0) AND_65 (c3540_wire_322, {c3540_wire_314, c3540_wire_323});
or_n #(2, 0, 0) OR_21 (c3540_wire_324, {c3540_wire_322, c3540_wire_310});
and_n #(2, 0, 0) AND_66 (c3540_wire_307, {c3540_wire_324, c3540_wire_325_0});
notg #(0, 0) NOT_129 (c3540_wire_312, c3540_wire_60_4);
notg #(0, 0) NOT_130 (c3540_wire_316, c3540_wire_120_2);
notg #(0, 0) NOT_131 (c3540_wire_323, c3540_wire_33_10);
notg #(0, 0) NOT_132 (c3540_wire_317, c3540_wire_18_3);
notg #(0, 0) NOT_133 (c3540_wire_319, c3540_wire_326_0);
notg #(0, 0) NOT_134 (c3540_wire_320, c3540_wire_325_1);
notg #(0, 0) NOT_135 (c3540_wire_321, c3540_wire_318_1);
notg #(0, 0) NOT_136 (c3540_wire_301, c3540_wire_327_0);
notg #(0, 0) NOT_137 (c3540_wire_328, c3540_wire_327_1);
or_n #(2, 0, 0) OR_22 (c3540_wire_304, {c3540_wire_327_2, c3540_wire_329});
and_n #(2, 0, 0) AND_67 (c3540_wire_327, {c3540_wire_330, c3540_wire_331});
and_n #(2, 0, 0) AND_68 (c3540_wire_332, {c3540_wire_333_0, c3540_wire_60_5});
or_n #(2, 0, 0) OR_23 (c3540_wire_334, {c3540_wire_332, c3540_wire_335});
and_n #(2, 0, 0) AND_69 (c3540_wire_336, {c3540_wire_54, c3540_wire_337});
or_n #(2, 0, 0) OR_24 (c3540_wire_338, {c3540_wire_336, c3540_wire_339});
or_n #(2, 0, 0) OR_25 (c3540_wire_330, {c3540_wire_338, c3540_wire_334});
and_n #(2, 0, 0) AND_70 (c3540_wire_335, {c3540_wire_340_0, c3540_wire_341_0});
notg #(0, 0) NOT_138 (c3540_wire_342, c3540_wire_341_1);
and_n #(2, 0, 0) AND_71 (c3540_wire_339, {c3540_wire_342, c3540_wire_9_3});
notg #(0, 0) NOT_139 (c3540_wire_343, c3540_wire_344_0);
and_n #(2, 0, 0) AND_72 (c3540_wire_55, {c3540_wire_343, c3540_wire_345});
notg #(0, 0) NOT_140 (c3540_wire_337, c3540_wire_60_6);
notg #(0, 0) NOT_141 (c3540_wire_331, c3540_wire_346_0);
and_n #(2, 0, 0) AND_73 (c3540_wire_347, {c3540_wire_298_0, c3540_wire_282});
or_n #(2, 0, 0) OR_26 (c3540_wire_348, {c3540_wire_298_1, c3540_wire_349_0});
bufg #(0, 0) BUF_9 (c3540_wire_350, G17_net_0);
notg #(0, 0) NOT_142 (c3540_wire_351, c3540_wire_352_0);
notg #(0, 0) NOT_143 (c3540_wire_353, c3540_wire_352_1);
or_n #(2, 0, 0) OR_27 (c3540_wire_354, {c3540_wire_352_2, c3540_wire_355});
and_n #(2, 0, 0) AND_74 (c3540_wire_352, {c3540_wire_356, c3540_wire_357});
and_n #(2, 0, 0) AND_75 (c3540_wire_358, {c3540_wire_9_4, c3540_wire_60_7});
or_n #(2, 0, 0) OR_28 (c3540_wire_359, {c3540_wire_358, c3540_wire_360});
and_n #(2, 0, 0) AND_76 (c3540_wire_361, {c3540_wire_102, c3540_wire_362});
or_n #(2, 0, 0) OR_29 (c3540_wire_363, {c3540_wire_361, c3540_wire_364});
or_n #(2, 0, 0) OR_30 (c3540_wire_356, {c3540_wire_363, c3540_wire_359});
and_n #(2, 0, 0) AND_77 (c3540_wire_360, {c3540_wire_340_1, c3540_wire_341_2});
notg #(0, 0) NOT_144 (c3540_wire_365, c3540_wire_341_3);
and_n #(2, 0, 0) AND_78 (c3540_wire_364, {c3540_wire_365, c3540_wire_10_2});
notg #(0, 0) NOT_145 (c3540_wire_366, c3540_wire_344_1);
and_n #(2, 0, 0) AND_79 (c3540_wire_103, {c3540_wire_366, c3540_wire_333_1});
notg #(0, 0) NOT_146 (c3540_wire_362, c3540_wire_60_8);
notg #(0, 0) NOT_147 (c3540_wire_357, c3540_wire_346_1);
and_n #(3, 0, 0) AND_80 (c3540_wire_367, {c3540_wire_73_1, c3540_wire_368, c3540_wire_369});
notg #(0, 0) NOT_148 (c3540_wire_370, c3540_wire_73_2);
and_n #(2, 0, 0) AND_81 (c3540_wire_371, {c3540_wire_73_3, c3540_wire_372});
or_n #(3, 0, 0) OR_31 (c3540_wire_73, {c3540_wire_373, c3540_wire_374, c3540_wire_375});
notg #(0, 0) NOT_149 (c3540_wire_376, c3540_wire_121_3);
and_n #(2, 0, 0) AND_82 (c3540_wire_377, {c3540_wire_376, c3540_wire_33_11});
and_n #(2, 0, 0) AND_83 (c3540_wire_378, {c3540_wire_379, c3540_wire_18_4});
or_n #(2, 0, 0) OR_32 (c3540_wire_380, {c3540_wire_378, c3540_wire_59});
and_n #(2, 0, 0) AND_84 (c3540_wire_373, {c3540_wire_381, c3540_wire_318_2});
and_n #(4, 0, 0) AND_85 (c3540_wire_374, {c3540_wire_382, c3540_wire_383, c3540_wire_384, c3540_wire_121_4});
and_n #(2, 0, 0) AND_86 (c3540_wire_385, {c3540_wire_380, c3540_wire_386});
or_n #(2, 0, 0) OR_33 (c3540_wire_387, {c3540_wire_385, c3540_wire_377});
and_n #(2, 0, 0) AND_87 (c3540_wire_375, {c3540_wire_387, c3540_wire_325_2});
notg #(0, 0) NOT_150 (c3540_wire_379, c3540_wire_60_9);
notg #(0, 0) NOT_151 (c3540_wire_386, c3540_wire_33_12);
notg #(0, 0) NOT_152 (c3540_wire_381, c3540_wire_121_5);
notg #(0, 0) NOT_153 (c3540_wire_382, c3540_wire_326_1);
notg #(0, 0) NOT_154 (c3540_wire_383, c3540_wire_325_3);
notg #(0, 0) NOT_155 (c3540_wire_384, c3540_wire_318_3);
notg #(0, 0) NOT_156 (c3540_wire_369, c3540_wire_388_0);
notg #(0, 0) NOT_157 (c3540_wire_389, c3540_wire_388_1);
or_n #(2, 0, 0) OR_34 (c3540_wire_372, {c3540_wire_388_2, c3540_wire_390});
and_n #(2, 0, 0) AND_88 (c3540_wire_388, {c3540_wire_391, c3540_wire_392});
and_n #(2, 0, 0) AND_89 (c3540_wire_393, {c3540_wire_10_3, c3540_wire_60_10});
or_n #(2, 0, 0) OR_35 (c3540_wire_394, {c3540_wire_393, c3540_wire_395});
and_n #(2, 0, 0) AND_90 (c3540_wire_396, {c3540_wire_127, c3540_wire_397});
or_n #(2, 0, 0) OR_36 (c3540_wire_398, {c3540_wire_396, c3540_wire_399});
or_n #(2, 0, 0) OR_37 (c3540_wire_391, {c3540_wire_398, c3540_wire_394});
and_n #(2, 0, 0) AND_91 (c3540_wire_395, {c3540_wire_340_2, c3540_wire_341_4});
notg #(0, 0) NOT_158 (c3540_wire_400, c3540_wire_341_5);
and_n #(2, 0, 0) AND_92 (c3540_wire_399, {c3540_wire_400, c3540_wire_401_0});
notg #(0, 0) NOT_159 (c3540_wire_402, c3540_wire_344_2);
and_n #(2, 0, 0) AND_93 (c3540_wire_128, {c3540_wire_402, c3540_wire_9_5});
notg #(0, 0) NOT_160 (c3540_wire_397, c3540_wire_60_11);
notg #(0, 0) NOT_161 (c3540_wire_392, c3540_wire_346_2);
and_n #(3, 0, 0) AND_94 (c3540_wire_403, {c3540_wire_75_1, c3540_wire_404, c3540_wire_405});
notg #(0, 0) NOT_162 (c3540_wire_406, c3540_wire_75_2);
and_n #(2, 0, 0) AND_95 (c3540_wire_407, {c3540_wire_75_3, c3540_wire_408});
or_n #(3, 0, 0) OR_38 (c3540_wire_75, {c3540_wire_409, c3540_wire_57, c3540_wire_410});
and_n #(2, 0, 0) AND_96 (c3540_wire_411, {c3540_wire_33_13, c3540_wire_325_4});
or_n #(2, 0, 0) OR_39 (c3540_wire_58, {c3540_wire_411, c3540_wire_412});
nor_n #(3, 0, 0) NOR_15 (c3540_wire_412, {c3540_wire_325_5, c3540_wire_326_2, c3540_wire_318_4});
and_n #(2, 0, 0) AND_97 (c3540_wire_409, {c3540_wire_56, c3540_wire_318_5});
and_n #(2, 0, 0) AND_98 (c3540_wire_413, {c3540_wire_104, c3540_wire_60_12});
or_n #(2, 0, 0) OR_40 (c3540_wire_414, {c3540_wire_413, c3540_wire_415});
nor_n #(2, 0, 0) NOR_16 (c3540_wire_415, {c3540_wire_60_13, c3540_wire_120_3});
and_n #(3, 0, 0) AND_99 (c3540_wire_410, {c3540_wire_414, c3540_wire_416, c3540_wire_325_6});
notg #(0, 0) NOT_163 (c3540_wire_416, c3540_wire_33_14);
notg #(0, 0) NOT_164 (c3540_wire_405, c3540_wire_417_0);
notg #(0, 0) NOT_165 (c3540_wire_418, c3540_wire_417_1);
or_n #(2, 0, 0) OR_41 (c3540_wire_408, {c3540_wire_417_2, c3540_wire_419});
and_n #(2, 0, 0) AND_100 (c3540_wire_417, {c3540_wire_420, c3540_wire_421});
and_n #(2, 0, 0) AND_101 (c3540_wire_422, {c3540_wire_401_1, c3540_wire_60_14});
or_n #(2, 0, 0) OR_42 (c3540_wire_423, {c3540_wire_422, c3540_wire_424});
and_n #(2, 0, 0) AND_102 (c3540_wire_425, {c3540_wire_183, c3540_wire_426});
or_n #(2, 0, 0) OR_43 (c3540_wire_427, {c3540_wire_425, c3540_wire_428});
or_n #(2, 0, 0) OR_44 (c3540_wire_420, {c3540_wire_427, c3540_wire_423});
and_n #(2, 0, 0) AND_103 (c3540_wire_424, {c3540_wire_340_3, c3540_wire_341_6});
notg #(0, 0) NOT_166 (c3540_wire_429, c3540_wire_341_7);
and_n #(2, 0, 0) AND_104 (c3540_wire_428, {c3540_wire_429, c3540_wire_430_0});
notg #(0, 0) NOT_167 (c3540_wire_431, c3540_wire_344_3);
and_n #(2, 0, 0) AND_105 (c3540_wire_184, {c3540_wire_431, c3540_wire_10_4});
notg #(0, 0) NOT_168 (c3540_wire_426, c3540_wire_60_15);
notg #(0, 0) NOT_169 (c3540_wire_421, c3540_wire_346_3);
and_n #(3, 0, 0) AND_106 (c3540_wire_432, {c3540_wire_69_1, c3540_wire_433, c3540_wire_434});
notg #(0, 0) NOT_170 (c3540_wire_435, c3540_wire_69_2);
and_n #(2, 0, 0) AND_107 (c3540_wire_436, {c3540_wire_69_3, c3540_wire_437});
or_n #(3, 0, 0) OR_45 (c3540_wire_69, {c3540_wire_438, c3540_wire_106, c3540_wire_439});
notg #(0, 0) NOT_171 (c3540_wire_440, c3540_wire_441);
and_n #(2, 0, 0) AND_108 (c3540_wire_442, {c3540_wire_440, c3540_wire_33_15});
or_n #(2, 0, 0) OR_46 (c3540_wire_443, {c3540_wire_442, c3540_wire_444});
and_n #(2, 0, 0) AND_109 (c3540_wire_445, {c3540_wire_129, c3540_wire_60_16});
or_n #(2, 0, 0) OR_47 (c3540_wire_446, {c3540_wire_445, c3540_wire_447});
nor_n #(2, 0, 0) NOR_17 (c3540_wire_447, {c3540_wire_60_17, c3540_wire_121_6});
and_n #(2, 0, 0) AND_110 (c3540_wire_438, {c3540_wire_105, c3540_wire_318_6});
and_n #(2, 0, 0) AND_111 (c3540_wire_444, {c3540_wire_446, c3540_wire_448});
and_n #(2, 0, 0) AND_112 (c3540_wire_439, {c3540_wire_443, c3540_wire_325_7});
notg #(0, 0) NOT_172 (c3540_wire_448, c3540_wire_33_16);
notg #(0, 0) NOT_173 (c3540_wire_107, c3540_wire_325_8);
notg #(0, 0) NOT_174 (c3540_wire_108, c3540_wire_449_0);
notg #(0, 0) NOT_175 (c3540_wire_109, c3540_wire_318_7);
notg #(0, 0) NOT_176 (c3540_wire_434, c3540_wire_450_0);
notg #(0, 0) NOT_177 (c3540_wire_451, c3540_wire_450_1);
or_n #(2, 0, 0) OR_48 (c3540_wire_437, {c3540_wire_450_2, c3540_wire_452});
and_n #(5, 0, 0) AND_113 (c3540_wire_453, {c3540_wire_450_3, c3540_wire_454_0, c3540_wire_455_0, c3540_wire_456_0, c3540_wire_150_4});
or_n #(2, 0, 0) OR_49 (c3540_wire_450, {c3540_wire_457, c3540_wire_458});
and_n #(2, 0, 0) AND_114 (c3540_wire_459, {c3540_wire_430_1, c3540_wire_60_18});
or_n #(2, 0, 0) OR_50 (c3540_wire_460, {c3540_wire_459, c3540_wire_461});
and_n #(3, 0, 0) AND_115 (c3540_wire_457, {c3540_wire_462, c3540_wire_463, c3540_wire_340_4});
or_n #(2, 0, 0) OR_51 (c3540_wire_464, {c3540_wire_460, c3540_wire_465});
and_n #(2, 0, 0) AND_116 (c3540_wire_465, {c3540_wire_206, c3540_wire_466});
and_n #(2, 0, 0) AND_117 (c3540_wire_458, {c3540_wire_464, c3540_wire_467});
or_n #(2, 0, 0) OR_52 (c3540_wire_468, {c3540_wire_1_4, c3540_wire_469_0});
and_n #(2, 0, 0) AND_118 (c3540_wire_461, {c3540_wire_468, c3540_wire_28_4});
notg #(0, 0) NOT_178 (c3540_wire_470, c3540_wire_344_4);
and_n #(2, 0, 0) AND_119 (c3540_wire_207, {c3540_wire_470, c3540_wire_401_2});
notg #(0, 0) NOT_179 (c3540_wire_466, c3540_wire_60_19);
notg #(0, 0) NOT_180 (c3540_wire_467, c3540_wire_346_4);
notg #(0, 0) NOT_181 (c3540_wire_462, c3540_wire_1_5);
notg #(0, 0) NOT_182 (c3540_wire_463, c3540_wire_469_1);
notg #(0, 0) NOT_183 (c3540_wire_471, c3540_wire_454_1);
notg #(0, 0) NOT_184 (c3540_wire_472, c3540_wire_454_2);
or_n #(2, 0, 0) OR_53 (c3540_wire_473, {c3540_wire_454_3, c3540_wire_474});
or_n #(2, 0, 0) OR_54 (c3540_wire_454, {c3540_wire_475, c3540_wire_476});
and_n #(2, 0, 0) AND_120 (c3540_wire_477, {c3540_wire_28_5, c3540_wire_60_20});
or_n #(2, 0, 0) OR_55 (c3540_wire_478, {c3540_wire_477, c3540_wire_479});
and_n #(2, 0, 0) AND_121 (c3540_wire_480, {c3540_wire_481, c3540_wire_430_2});
or_n #(2, 0, 0) OR_56 (c3540_wire_482, {c3540_wire_480, c3540_wire_483_0});
and_n #(4, 0, 0) AND_122 (c3540_wire_475, {c3540_wire_484, c3540_wire_485, c3540_wire_486, c3540_wire_340_5});
or_n #(2, 0, 0) OR_57 (c3540_wire_487, {c3540_wire_478, c3540_wire_488});
and_n #(2, 0, 0) AND_123 (c3540_wire_488, {c3540_wire_482, c3540_wire_489});
and_n #(2, 0, 0) AND_124 (c3540_wire_476, {c3540_wire_487, c3540_wire_490});
notg #(0, 0) NOT_185 (c3540_wire_491, c3540_wire_492_0);
and_n #(2, 0, 0) AND_125 (c3540_wire_479, {c3540_wire_491, c3540_wire_111_2});
notg #(0, 0) NOT_186 (c3540_wire_481, c3540_wire_344_5);
notg #(0, 0) NOT_187 (c3540_wire_489, c3540_wire_60_21);
notg #(0, 0) NOT_188 (c3540_wire_490, c3540_wire_346_5);
notg #(0, 0) NOT_189 (c3540_wire_484, c3540_wire_1_6);
notg #(0, 0) NOT_190 (c3540_wire_485, c3540_wire_38_1);
notg #(0, 0) NOT_191 (c3540_wire_486, c3540_wire_469_2);
and_n #(3, 0, 0) AND_126 (c3540_wire_493, {c3540_wire_79_1, c3540_wire_494, c3540_wire_495});
notg #(0, 0) NOT_192 (c3540_wire_496, c3540_wire_79_2);
and_n #(2, 0, 0) AND_127 (c3540_wire_497, {c3540_wire_79_3, c3540_wire_498});
or_n #(3, 0, 0) OR_58 (c3540_wire_79, {c3540_wire_186, c3540_wire_499, c3540_wire_500});
and_n #(2, 0, 0) AND_128 (c3540_wire_501, {c3540_wire_33_17, c3540_wire_325_9});
or_n #(2, 0, 0) OR_59 (c3540_wire_502, {c3540_wire_501, c3540_wire_318_8});
and_n #(2, 0, 0) AND_129 (c3540_wire_499, {c3540_wire_502, c3540_wire_185});
nor_n #(2, 0, 0) NOR_18 (c3540_wire_503, {c3540_wire_5_10, c3540_wire_60_22});
or_n #(2, 0, 0) OR_60 (c3540_wire_504, {c3540_wire_503, c3540_wire_211});
and_n #(3, 0, 0) AND_130 (c3540_wire_500, {c3540_wire_504, c3540_wire_505, c3540_wire_325_10});
notg #(0, 0) NOT_193 (c3540_wire_505, c3540_wire_33_18);
notg #(0, 0) NOT_194 (c3540_wire_187, c3540_wire_325_11);
notg #(0, 0) NOT_195 (c3540_wire_188, c3540_wire_449_1);
notg #(0, 0) NOT_196 (c3540_wire_189, c3540_wire_318_9);
notg #(0, 0) NOT_197 (c3540_wire_495, c3540_wire_455_1);
notg #(0, 0) NOT_198 (c3540_wire_506, c3540_wire_455_2);
or_n #(2, 0, 0) OR_61 (c3540_wire_498, {c3540_wire_455_3, c3540_wire_507});
or_n #(2, 0, 0) OR_62 (c3540_wire_455, {c3540_wire_508, c3540_wire_509});
and_n #(2, 0, 0) AND_131 (c3540_wire_510, {c3540_wire_111_3, c3540_wire_60_23});
or_n #(2, 0, 0) OR_63 (c3540_wire_511, {c3540_wire_510, c3540_wire_512});
and_n #(2, 0, 0) AND_132 (c3540_wire_513, {c3540_wire_514, c3540_wire_28_6});
or_n #(2, 0, 0) OR_64 (c3540_wire_515, {c3540_wire_513, c3540_wire_516_0});
and_n #(4, 0, 0) AND_133 (c3540_wire_508, {c3540_wire_517, c3540_wire_518, c3540_wire_519, c3540_wire_340_6});
or_n #(2, 0, 0) OR_65 (c3540_wire_520, {c3540_wire_511, c3540_wire_521});
and_n #(2, 0, 0) AND_134 (c3540_wire_521, {c3540_wire_515, c3540_wire_522});
and_n #(2, 0, 0) AND_135 (c3540_wire_509, {c3540_wire_520, c3540_wire_523});
notg #(0, 0) NOT_199 (c3540_wire_524, c3540_wire_492_1);
and_n #(2, 0, 0) AND_136 (c3540_wire_512, {c3540_wire_524, c3540_wire_115_2});
notg #(0, 0) NOT_200 (c3540_wire_514, c3540_wire_344_6);
notg #(0, 0) NOT_201 (c3540_wire_522, c3540_wire_60_24);
notg #(0, 0) NOT_202 (c3540_wire_523, c3540_wire_346_6);
notg #(0, 0) NOT_203 (c3540_wire_517, c3540_wire_1_7);
notg #(0, 0) NOT_204 (c3540_wire_518, c3540_wire_38_2);
notg #(0, 0) NOT_205 (c3540_wire_519, c3540_wire_469_3);
and_n #(3, 0, 0) AND_137 (c3540_wire_525, {c3540_wire_71_1, c3540_wire_526, c3540_wire_527});
notg #(0, 0) NOT_206 (c3540_wire_528, c3540_wire_71_2);
and_n #(2, 0, 0) AND_138 (c3540_wire_529, {c3540_wire_71_3, c3540_wire_530});
or_n #(3, 0, 0) OR_66 (c3540_wire_71, {c3540_wire_531, c3540_wire_209, c3540_wire_532});
and_n #(2, 0, 0) AND_139 (c3540_wire_533, {c3540_wire_33_19, c3540_wire_325_12});
or_n #(2, 0, 0) OR_67 (c3540_wire_210, {c3540_wire_533, c3540_wire_534});
nor_n #(3, 0, 0) NOR_19 (c3540_wire_534, {c3540_wire_449_2, c3540_wire_325_13, c3540_wire_318_10});
and_n #(2, 0, 0) AND_140 (c3540_wire_531, {c3540_wire_208, c3540_wire_318_11});
nor_n #(2, 0, 0) NOR_20 (c3540_wire_535, {c3540_wire_99_11, c3540_wire_60_25});
or_n #(2, 0, 0) OR_68 (c3540_wire_536, {c3540_wire_535, c3540_wire_537});
and_n #(3, 0, 0) AND_141 (c3540_wire_532, {c3540_wire_536, c3540_wire_538, c3540_wire_325_14});
and_n #(2, 0, 0) AND_142 (c3540_wire_537, {c3540_wire_483_1, c3540_wire_60_26});
notg #(0, 0) NOT_207 (c3540_wire_538, c3540_wire_33_20);
notg #(0, 0) NOT_208 (c3540_wire_527, c3540_wire_456_1);
notg #(0, 0) NOT_209 (c3540_wire_539, c3540_wire_456_2);
or_n #(2, 0, 0) OR_69 (c3540_wire_530, {c3540_wire_456_3, c3540_wire_540});
or_n #(2, 0, 0) OR_70 (c3540_wire_456, {c3540_wire_541, c3540_wire_542});
and_n #(2, 0, 0) AND_143 (c3540_wire_543, {c3540_wire_115_3, c3540_wire_60_27});
or_n #(2, 0, 0) OR_71 (c3540_wire_544, {c3540_wire_543, c3540_wire_545});
and_n #(2, 0, 0) AND_144 (c3540_wire_546, {c3540_wire_547, c3540_wire_111_4});
or_n #(2, 0, 0) OR_72 (c3540_wire_548, {c3540_wire_546, c3540_wire_549_0});
and_n #(4, 0, 0) AND_145 (c3540_wire_541, {c3540_wire_550, c3540_wire_551, c3540_wire_552, c3540_wire_340_7});
or_n #(2, 0, 0) OR_73 (c3540_wire_553, {c3540_wire_544, c3540_wire_554});
and_n #(2, 0, 0) AND_146 (c3540_wire_554, {c3540_wire_548, c3540_wire_555});
and_n #(2, 0, 0) AND_147 (c3540_wire_542, {c3540_wire_553, c3540_wire_556});
notg #(0, 0) NOT_210 (c3540_wire_557, c3540_wire_492_2);
and_n #(2, 0, 0) AND_148 (c3540_wire_545, {c3540_wire_557, c3540_wire_116_2});
notg #(0, 0) NOT_211 (c3540_wire_547, c3540_wire_344_7);
notg #(0, 0) NOT_212 (c3540_wire_555, c3540_wire_60_28);
notg #(0, 0) NOT_213 (c3540_wire_556, c3540_wire_346_7);
notg #(0, 0) NOT_214 (c3540_wire_550, c3540_wire_1_8);
notg #(0, 0) NOT_215 (c3540_wire_551, c3540_wire_38_3);
notg #(0, 0) NOT_216 (c3540_wire_552, c3540_wire_469_4);
notg #(0, 0) NOT_217 (c3540_wire_558, c3540_wire_559);
or_n #(3, 0, 0) OR_74 (c3540_wire_559, {c3540_wire_560, c3540_wire_561, c3540_wire_146});
and_n #(2, 0, 0) AND_149 (c3540_wire_561, {c3540_wire_43, c3540_wire_562});
nor_n #(3, 0, 0) NOR_21 (c3540_wire_560, {c3540_wire_39_5, c3540_wire_13, c3540_wire_30_1});
or_n #(2, 0, 0) OR_75 (c3540_wire_562, {c3540_wire_111_5, c3540_wire_115_4});
notg #(0, 0) NOT_218 (c3540_wire_147, c3540_wire_18_5);
and_n #(2, 0, 0) AND_150 (c3540_wire_563, {c3540_wire_350_0, c3540_wire_270});
and_n #(2, 0, 0) AND_151 (c3540_wire_564, {c3540_wire_350_1, c3540_wire_283});
or_n #(2, 0, 0) OR_76 (c3540_wire_565, {c3540_wire_350_2, c3540_wire_313_1});
bufg #(0, 0) BUF_10 (c3540_wire_566, G18_net_0);
or_n #(2, 0, 0) OR_77 (c3540_wire_53, {c3540_wire_216, c3540_wire_567});
nor_n #(2, 0, 0) NOR_22 (c3540_wire_567, {c3540_wire_215_2, c3540_wire_121_7});
or_n #(2, 0, 0) OR_78 (c3540_wire_568, {c3540_wire_217, c3540_wire_569});
or_n #(2, 0, 0) OR_79 (c3540_wire_221, {c3540_wire_52, c3540_wire_570});
nor_n #(2, 0, 0) NOR_23 (c3540_wire_570, {c3540_wire_568, c3540_wire_2_12});
nor_n #(2, 0, 0) NOR_24 (c3540_wire_569, {c3540_wire_215_3, c3540_wire_121_8});
or_n #(2, 0, 0) OR_80 (c3540_wire_571, {c3540_wire_566_0, c3540_wire_572_0});
and_n #(2, 0, 0) AND_152 (c3540_wire_573, {c3540_wire_566_1, c3540_wire_271});
or_n #(2, 0, 0) OR_81 (c3540_wire_574, {c3540_wire_566_2, c3540_wire_572_1});
and_n #(2, 0, 0) AND_153 (c3540_wire_575, {c3540_wire_566_3, c3540_wire_285});
bufg #(0, 0) BUF_11 (c3540_wire_297, G19_net_0);
or_n #(2, 0, 0) OR_82 (c3540_wire_576, {c3540_wire_297_1, c3540_wire_577});
and_n #(2, 0, 0) AND_154 (c3540_wire_578, {c3540_wire_297_2, c3540_wire_284});
and_n #(2, 0, 0) AND_155 (c3540_wire_579, {c3540_wire_297_3, c3540_wire_273});
or_n #(2, 0, 0) OR_83 (c3540_wire_580, {c3540_wire_297_4, c3540_wire_581});
notg #(0, 0) NOT_219 (c3540_wire_582, c3540_wire_1_9);
notg #(0, 0) NOT_220 (c3540_wire_583, c3540_wire_1_10);
and_n #(2, 0, 0) AND_156 (c3540_wire_325, {c3540_wire_1_11, c3540_wire_584});
notg #(0, 0) NOT_221 (c3540_wire_585, c3540_wire_1_12);
notg #(0, 0) NOT_222 (c3540_wire_586, c3540_wire_1_13);
and_n #(2, 0, 0) AND_157 (c3540_wire_587, {c3540_wire_1_14, c3540_wire_32_4});
notg #(0, 0) NOT_223 (c3540_wire_588, c3540_wire_1_15);
notg #(0, 0) NOT_224 (c3540_wire_589, c3540_wire_1_16);
notg #(0, 0) NOT_225 (c3540_wire_590, c3540_wire_1_17);
notg #(0, 0) NOT_226 (c3540_wire_591, c3540_wire_1_18);
notg #(0, 0) NOT_227 (c3540_wire_592, c3540_wire_1_19);
notg #(0, 0) NOT_228 (c3540_wire_593, c3540_wire_1_20);
or_n #(2, 0, 0) OR_84 (c3540_wire_594, {c3540_wire_1_21, c3540_wire_595});
bufg #(0, 0) BUF_12 (c3540_wire_32, G2_net_0);
bufg #(0, 0) BUF_13 (c3540_wire_349, G20_net_0);
xor_n #(2, 0, 0) XOR_5 (c3540_wire_596, {c3540_wire_44, c3540_wire_597_0});
or_n #(2, 0, 0) OR_85 (c3540_wire_138, {c3540_wire_196, c3540_wire_598});
and_n #(2, 0, 0) AND_158 (c3540_wire_599, {c3540_wire_401_3, c3540_wire_430_3});
or_n #(2, 0, 0) OR_86 (c3540_wire_197, {c3540_wire_599, c3540_wire_600});
or_n #(2, 0, 0) OR_87 (c3540_wire_601, {c3540_wire_602, c3540_wire_603});
nor_n #(2, 0, 0) NOR_25 (c3540_wire_598, {c3540_wire_601, c3540_wire_11_1});
nor_n #(2, 0, 0) NOR_26 (c3540_wire_600, {c3540_wire_401_4, c3540_wire_430_4});
and_n #(2, 0, 0) AND_159 (c3540_wire_602, {c3540_wire_401_5, c3540_wire_430_5});
nor_n #(2, 0, 0) NOR_27 (c3540_wire_603, {c3540_wire_401_6, c3540_wire_430_6});
and_n #(2, 0, 0) AND_160 (c3540_wire_604, {c3540_wire_349_1, c3540_wire_264});
and_n #(2, 0, 0) AND_161 (c3540_wire_605, {c3540_wire_349_2, c3540_wire_272});
or_n #(2, 0, 0) OR_88 (c3540_wire_606, {c3540_wire_349_3, c3540_wire_607});
and_n #(2, 0, 0) AND_162 (c3540_wire_608, {c3540_wire_349_4, c3540_wire_289});
or_n #(2, 0, 0) OR_89 (c3540_wire_609, {c3540_wire_349_5, c3540_wire_610});
bufg #(0, 0) BUF_14 (c3540_wire_313, G21_net_0);
or_n #(6, 0, 0) OR_90 (c3540_wire_611, {c3540_wire_347, c3540_wire_604, c3540_wire_612, c3540_wire_613, c3540_wire_614, c3540_wire_563});
notg #(0, 0) NOT_229 (c3540_wire_615, c3540_wire_611);
and_n #(2, 0, 0) AND_163 (c3540_wire_612, {c3540_wire_262, c3540_wire_313_2});
and_n #(2, 0, 0) AND_164 (c3540_wire_613, {c3540_wire_296, c3540_wire_223});
and_n #(2, 0, 0) AND_165 (c3540_wire_614, {c3540_wire_571, c3540_wire_245});
or_n #(2, 0, 0) OR_91 (c3540_wire_616, {c3540_wire_617, c3540_wire_618});
or_n #(4, 0, 0) OR_92 (c3540_wire_617, {c3540_wire_564, c3540_wire_619, c3540_wire_620, c3540_wire_573});
and_n #(2, 0, 0) AND_166 (c3540_wire_619, {c3540_wire_265, c3540_wire_313_3});
and_n #(2, 0, 0) AND_167 (c3540_wire_620, {c3540_wire_263, c3540_wire_572_2});
and_n #(2, 0, 0) AND_168 (c3540_wire_621, {c3540_wire_348, c3540_wire_225});
or_n #(2, 0, 0) OR_93 (c3540_wire_618, {c3540_wire_621, c3540_wire_622});
and_n #(2, 0, 0) AND_169 (c3540_wire_622, {c3540_wire_576, c3540_wire_246});
notg #(0, 0) NOT_230 (c3540_wire_577, c3540_wire_18_6);
or_n #(2, 0, 0) OR_94 (c3540_wire_623, {c3540_wire_624, c3540_wire_625});
or_n #(4, 0, 0) OR_95 (c3540_wire_624, {c3540_wire_579, c3540_wire_575, c3540_wire_626, c3540_wire_627});
and_n #(2, 0, 0) AND_170 (c3540_wire_626, {c3540_wire_266, c3540_wire_572_3});
and_n #(2, 0, 0) AND_171 (c3540_wire_627, {c3540_wire_565, c3540_wire_227});
and_n #(2, 0, 0) AND_172 (c3540_wire_628, {c3540_wire_606, c3540_wire_248});
nor_n #(2, 0, 0) NOR_28 (c3540_wire_629, {c3540_wire_153_2, c3540_wire_18_7});
or_n #(2, 0, 0) OR_96 (c3540_wire_625, {c3540_wire_629, c3540_wire_628});
notg #(0, 0) NOT_231 (c3540_wire_607, c3540_wire_120_4);
or_n #(3, 0, 0) OR_97 (c3540_wire_630, {c3540_wire_631, c3540_wire_632, c3540_wire_633});
nor_n #(2, 0, 0) NOR_29 (c3540_wire_634, {c3540_wire_120_5, c3540_wire_153_3});
or_n #(2, 0, 0) OR_98 (c3540_wire_631, {c3540_wire_605, c3540_wire_578});
and_n #(2, 0, 0) AND_173 (c3540_wire_635, {c3540_wire_574, c3540_wire_226});
or_n #(2, 0, 0) OR_99 (c3540_wire_633, {c3540_wire_635, c3540_wire_636});
or_n #(2, 0, 0) OR_100 (c3540_wire_637, {c3540_wire_638, c3540_wire_313_4});
and_n #(2, 0, 0) AND_174 (c3540_wire_636, {c3540_wire_637, c3540_wire_247});
nor_n #(2, 0, 0) NOR_30 (c3540_wire_639, {c3540_wire_155_6, c3540_wire_18_8});
or_n #(2, 0, 0) OR_101 (c3540_wire_632, {c3540_wire_639, c3540_wire_634});
notg #(0, 0) NOT_232 (c3540_wire_638, c3540_wire_121_9);
or_n #(2, 0, 0) OR_102 (c3540_wire_640, {c3540_wire_641, c3540_wire_642});
or_n #(2, 0, 0) OR_103 (c3540_wire_643, {c3540_wire_100, c3540_wire_483_2});
nor_n #(2, 0, 0) NOR_31 (c3540_wire_644, {c3540_wire_153_4, c3540_wire_121_10});
nor_n #(2, 0, 0) NOR_32 (c3540_wire_645, {c3540_wire_181_10, c3540_wire_161_14});
and_n #(2, 0, 0) AND_175 (c3540_wire_646, {c3540_wire_643, c3540_wire_229});
nand_n #(2, 0, 0) NAND_1 (c3540_wire_647, {c3540_wire_99_12, c3540_wire_120_6});
and_n #(2, 0, 0) AND_176 (c3540_wire_648, {c3540_wire_647, c3540_wire_250});
nor_n #(2, 0, 0) NOR_33 (c3540_wire_649, {c3540_wire_2_13, c3540_wire_155_7});
or_n #(2, 0, 0) OR_104 (c3540_wire_650, {c3540_wire_649, c3540_wire_651});
nor_n #(2, 0, 0) NOR_34 (c3540_wire_651, {c3540_wire_123_11, c3540_wire_157_12});
or_n #(2, 0, 0) OR_105 (c3540_wire_641, {c3540_wire_644, c3540_wire_645});
or_n #(3, 0, 0) OR_106 (c3540_wire_642, {c3540_wire_646, c3540_wire_648, c3540_wire_650});
or_n #(5, 0, 0) OR_107 (c3540_wire_652, {c3540_wire_653, c3540_wire_654, c3540_wire_655, c3540_wire_656, c3540_wire_657});
notg #(0, 0) NOT_233 (c3540_wire_658, c3540_wire_652);
and_n #(2, 0, 0) AND_177 (c3540_wire_653, {c3540_wire_288, c3540_wire_483_3});
nor_n #(2, 0, 0) NOR_35 (c3540_wire_659, {c3540_wire_157_13, c3540_wire_181_11});
nor_n #(2, 0, 0) NOR_36 (c3540_wire_660, {c3540_wire_5_11, c3540_wire_155_8});
or_n #(2, 0, 0) OR_108 (c3540_wire_661, {c3540_wire_126, c3540_wire_516_1});
and_n #(2, 0, 0) AND_178 (c3540_wire_655, {c3540_wire_661, c3540_wire_231});
nand_n #(2, 0, 0) NAND_2 (c3540_wire_662, {c3540_wire_123_12, c3540_wire_121_11});
and_n #(2, 0, 0) AND_179 (c3540_wire_656, {c3540_wire_662, c3540_wire_252});
nor_n #(2, 0, 0) NOR_37 (c3540_wire_654, {c3540_wire_2_14, c3540_wire_153_5});
or_n #(2, 0, 0) OR_109 (c3540_wire_657, {c3540_wire_659, c3540_wire_660});
or_n #(3, 0, 0) OR_110 (c3540_wire_663, {c3540_wire_664, c3540_wire_665, c3540_wire_666});
notg #(0, 0) NOT_234 (c3540_wire_667, c3540_wire_663);
and_n #(2, 0, 0) AND_180 (c3540_wire_668, {c3540_wire_286, c3540_wire_516_2});
nor_n #(2, 0, 0) NOR_38 (c3540_wire_669, {c3540_wire_5_12, c3540_wire_153_6});
or_n #(2, 0, 0) OR_111 (c3540_wire_664, {c3540_wire_668, c3540_wire_670});
and_n #(2, 0, 0) AND_181 (c3540_wire_670, {c3540_wire_274, c3540_wire_483_4});
or_n #(2, 0, 0) OR_112 (c3540_wire_671, {c3540_wire_182, c3540_wire_549_1});
and_n #(2, 0, 0) AND_182 (c3540_wire_672, {c3540_wire_671, c3540_wire_228});
nand_n #(2, 0, 0) NAND_3 (c3540_wire_673, {c3540_wire_2_15, c3540_wire_181_12});
and_n #(2, 0, 0) AND_183 (c3540_wire_674, {c3540_wire_673, c3540_wire_249});
nor_n #(2, 0, 0) NOR_39 (c3540_wire_675, {c3540_wire_99_13, c3540_wire_155_9});
or_n #(2, 0, 0) OR_113 (c3540_wire_665, {c3540_wire_675, c3540_wire_669});
or_n #(2, 0, 0) OR_114 (c3540_wire_666, {c3540_wire_672, c3540_wire_674});
or_n #(3, 0, 0) OR_115 (c3540_wire_676, {c3540_wire_677, c3540_wire_678, c3540_wire_679});
notg #(0, 0) NOT_235 (c3540_wire_680, c3540_wire_676);
and_n #(2, 0, 0) AND_184 (c3540_wire_681, {c3540_wire_287, c3540_wire_549_2});
nor_n #(2, 0, 0) NOR_40 (c3540_wire_682, {c3540_wire_153_7, c3540_wire_99_14});
or_n #(2, 0, 0) OR_116 (c3540_wire_677, {c3540_wire_681, c3540_wire_683});
and_n #(2, 0, 0) AND_185 (c3540_wire_683, {c3540_wire_275, c3540_wire_516_3});
or_n #(2, 0, 0) OR_117 (c3540_wire_684, {c3540_wire_205, c3540_wire_685_0});
and_n #(2, 0, 0) AND_186 (c3540_wire_686, {c3540_wire_684, c3540_wire_230});
or_n #(2, 0, 0) OR_118 (c3540_wire_687, {c3540_wire_101, c3540_wire_483_5});
and_n #(2, 0, 0) AND_187 (c3540_wire_688, {c3540_wire_687, c3540_wire_251});
nor_n #(2, 0, 0) NOR_41 (c3540_wire_689, {c3540_wire_123_13, c3540_wire_155_10});
or_n #(2, 0, 0) OR_119 (c3540_wire_678, {c3540_wire_689, c3540_wire_682});
or_n #(2, 0, 0) OR_120 (c3540_wire_679, {c3540_wire_686, c3540_wire_688});
and_n #(2, 0, 0) AND_188 (c3540_wire_690, {c3540_wire_313_5, c3540_wire_276});
and_n #(2, 0, 0) AND_189 (c3540_wire_691, {c3540_wire_313_6, c3540_wire_291});
or_n #(2, 0, 0) OR_121 (c3540_wire_692, {c3540_wire_313_7, c3540_wire_693});
bufg #(0, 0) BUF_15 (c3540_wire_572, G22_net_0);
and_n #(3, 0, 0) AND_190 (c3540_wire_694, {c3540_wire_47_1, c3540_wire_695, c3540_wire_351});
notg #(0, 0) NOT_236 (c3540_wire_696, c3540_wire_47_2);
and_n #(2, 0, 0) AND_191 (c3540_wire_697, {c3540_wire_47_3, c3540_wire_354});
or_n #(3, 0, 0) OR_122 (c3540_wire_47, {c3540_wire_698, c3540_wire_699, c3540_wire_700});
xor_n #(2, 0, 0) XOR_6 (c3540_wire_701, {c3540_wire_120_7, c3540_wire_121_12});
and_n #(2, 0, 0) AND_192 (c3540_wire_702, {c3540_wire_701, c3540_wire_33_21});
and_n #(2, 0, 0) AND_193 (c3540_wire_703, {c3540_wire_704, c3540_wire_572_4});
or_n #(2, 0, 0) OR_123 (c3540_wire_705, {c3540_wire_703, c3540_wire_706});
and_n #(2, 0, 0) AND_194 (c3540_wire_706, {c3540_wire_707, c3540_wire_60_29});
and_n #(2, 0, 0) AND_195 (c3540_wire_698, {c3540_wire_708, c3540_wire_318_12});
and_n #(4, 0, 0) AND_196 (c3540_wire_699, {c3540_wire_709, c3540_wire_710, c3540_wire_711, c3540_wire_120_8});
and_n #(2, 0, 0) AND_197 (c3540_wire_712, {c3540_wire_705, c3540_wire_713});
or_n #(2, 0, 0) OR_124 (c3540_wire_714, {c3540_wire_712, c3540_wire_702});
and_n #(2, 0, 0) AND_198 (c3540_wire_700, {c3540_wire_714, c3540_wire_325_15});
notg #(0, 0) NOT_237 (c3540_wire_704, c3540_wire_60_30);
notg #(0, 0) NOT_238 (c3540_wire_707, c3540_wire_121_13);
notg #(0, 0) NOT_239 (c3540_wire_713, c3540_wire_33_22);
notg #(0, 0) NOT_240 (c3540_wire_708, c3540_wire_120_9);
notg #(0, 0) NOT_241 (c3540_wire_709, c3540_wire_326_3);
notg #(0, 0) NOT_242 (c3540_wire_710, c3540_wire_325_16);
notg #(0, 0) NOT_243 (c3540_wire_711, c3540_wire_318_13);
and_n #(3, 0, 0) AND_199 (c3540_wire_715, {c3540_wire_77_1, c3540_wire_716, c3540_wire_471});
notg #(0, 0) NOT_244 (c3540_wire_717, c3540_wire_77_2);
and_n #(2, 0, 0) AND_200 (c3540_wire_718, {c3540_wire_77_3, c3540_wire_473});
or_n #(3, 0, 0) OR_125 (c3540_wire_77, {c3540_wire_719, c3540_wire_131, c3540_wire_720});
or_n #(2, 0, 0) OR_126 (c3540_wire_721, {c3540_wire_202, c3540_wire_722});
and_n #(2, 0, 0) AND_201 (c3540_wire_719, {c3540_wire_130, c3540_wire_318_14});
or_n #(2, 0, 0) OR_127 (c3540_wire_723, {c3540_wire_190, c3540_wire_61});
and_n #(2, 0, 0) AND_202 (c3540_wire_722, {c3540_wire_723, c3540_wire_724});
and_n #(2, 0, 0) AND_203 (c3540_wire_720, {c3540_wire_721, c3540_wire_325_17});
notg #(0, 0) NOT_245 (c3540_wire_62, c3540_wire_60_31);
notg #(0, 0) NOT_246 (c3540_wire_724, c3540_wire_33_23);
notg #(0, 0) NOT_247 (c3540_wire_132, c3540_wire_325_18);
notg #(0, 0) NOT_248 (c3540_wire_133, c3540_wire_449_3);
notg #(0, 0) NOT_249 (c3540_wire_134, c3540_wire_318_15);
or_n #(2, 0, 0) OR_128 (c3540_wire_725, {c3540_wire_572_5, c3540_wire_64});
and_n #(2, 0, 0) AND_204 (c3540_wire_726, {c3540_wire_572_6, c3540_wire_278});
and_n #(2, 0, 0) AND_205 (c3540_wire_727, {c3540_wire_572_7, c3540_wire_293});
or_n #(2, 0, 0) OR_129 (c3540_wire_728, {c3540_wire_572_8, c3540_wire_65});
bufg #(0, 0) BUF_16 (c3540_wire_178, G23_net_0);
notg #(0, 0) NOT_250 (c3540_wire_729, c3540_wire_299);
or_n #(2, 0, 0) OR_130 (c3540_wire_300, {c3540_wire_178_1, c3540_wire_150_5});
notg #(0, 0) NOT_251 (c3540_wire_730, c3540_wire_367_0);
notg #(0, 0) NOT_252 (c3540_wire_88, c3540_wire_367_1);
and_n #(2, 0, 0) AND_206 (c3540_wire_731, {c3540_wire_367_2, c3540_wire_732_0});
or_n #(2, 0, 0) OR_131 (c3540_wire_368, {c3540_wire_178_2, c3540_wire_150_6});
and_n #(2, 0, 0) AND_207 (c3540_wire_733, {c3540_wire_403_0, c3540_wire_66});
or_n #(2, 0, 0) OR_132 (c3540_wire_404, {c3540_wire_178_3, c3540_wire_150_7});
notg #(0, 0) NOT_253 (c3540_wire_734, c3540_wire_432);
or_n #(2, 0, 0) OR_133 (c3540_wire_433, {c3540_wire_178_4, c3540_wire_150_8});
notg #(0, 0) NOT_254 (c3540_wire_735, c3540_wire_493_0);
and_n #(2, 0, 0) AND_208 (c3540_wire_736, {c3540_wire_493_1, c3540_wire_90});
notg #(0, 0) NOT_255 (c3540_wire_737, c3540_wire_493_2);
or_n #(2, 0, 0) OR_134 (c3540_wire_494, {c3540_wire_178_5, c3540_wire_150_9});
and_n #(2, 0, 0) AND_209 (c3540_wire_738, {c3540_wire_525_0, c3540_wire_67});
and_n #(2, 0, 0) AND_210 (c3540_wire_739, {c3540_wire_525_1, c3540_wire_83_1});
or_n #(2, 0, 0) OR_135 (c3540_wire_526, {c3540_wire_178_6, c3540_wire_150_10});
xor_n #(2, 0, 0) XOR_7 (c3540_wire_732, {c3540_wire_46, c3540_wire_740_0});
or_n #(2, 0, 0) OR_136 (c3540_wire_716, {c3540_wire_178_7, c3540_wire_150_11});
or_n #(2, 0, 0) OR_137 (c3540_wire_695, {c3540_wire_178_8, c3540_wire_150_12});
bufg #(0, 0) BUF_17 (c3540_wire_150, G24_net_0);
and_n #(4, 0, 0) AND_211 (c3540_wire_741, {c3540_wire_597_1, c3540_wire_742_0, c3540_wire_743_0, c3540_wire_740_1});
or_n #(2, 0, 0) OR_138 (c3540_wire_597, {c3540_wire_744, c3540_wire_303});
notg #(0, 0) NOT_256 (c3540_wire_745, c3540_wire_597_2);
nor_n #(2, 0, 0) NOR_42 (c3540_wire_329, {c3540_wire_178_9, c3540_wire_150_13});
or_n #(2, 0, 0) OR_139 (c3540_wire_746, {c3540_wire_149_4, c3540_wire_151_6});
and_n #(3, 0, 0) AND_212 (c3540_wire_744, {c3540_wire_746, c3540_wire_328, c3540_wire_302});
or_n #(2, 0, 0) OR_140 (c3540_wire_742, {c3540_wire_747, c3540_wire_371});
notg #(0, 0) NOT_257 (c3540_wire_748, c3540_wire_742_1);
and_n #(2, 0, 0) AND_213 (c3540_wire_749, {c3540_wire_742_2, c3540_wire_750});
nor_n #(2, 0, 0) NOR_43 (c3540_wire_390, {c3540_wire_178_10, c3540_wire_150_14});
or_n #(2, 0, 0) OR_141 (c3540_wire_751, {c3540_wire_149_5, c3540_wire_151_7});
and_n #(3, 0, 0) AND_214 (c3540_wire_747, {c3540_wire_751, c3540_wire_389, c3540_wire_370});
or_n #(2, 0, 0) OR_142 (c3540_wire_743, {c3540_wire_752, c3540_wire_407});
notg #(0, 0) NOT_258 (c3540_wire_753, c3540_wire_743_1);
and_n #(2, 0, 0) AND_215 (c3540_wire_754, {c3540_wire_743_2, c3540_wire_755});
nor_n #(2, 0, 0) NOR_44 (c3540_wire_419, {c3540_wire_178_11, c3540_wire_150_15});
or_n #(2, 0, 0) OR_143 (c3540_wire_756, {c3540_wire_149_6, c3540_wire_151_8});
and_n #(3, 0, 0) AND_216 (c3540_wire_752, {c3540_wire_756, c3540_wire_418, c3540_wire_406});
or_n #(2, 0, 0) OR_144 (c3540_wire_82, {c3540_wire_757, c3540_wire_436});
and_n #(5, 0, 0) AND_217 (c3540_wire_758, {c3540_wire_82_1, c3540_wire_83_2, c3540_wire_84_1, c3540_wire_85_1, c3540_wire_741_0});
notg #(0, 0) NOT_259 (c3540_wire_759, c3540_wire_82_2);
and_n #(2, 0, 0) AND_218 (c3540_wire_760, {c3540_wire_82_3, c3540_wire_761});
notg #(0, 0) NOT_260 (c3540_wire_762, c3540_wire_82_4);
nor_n #(2, 0, 0) NOR_45 (c3540_wire_452, {c3540_wire_178_12, c3540_wire_150_16});
or_n #(2, 0, 0) OR_145 (c3540_wire_763, {c3540_wire_149_7, c3540_wire_151_9});
and_n #(3, 0, 0) AND_219 (c3540_wire_757, {c3540_wire_763, c3540_wire_451, c3540_wire_435});
or_n #(2, 0, 0) OR_146 (c3540_wire_83, {c3540_wire_764, c3540_wire_497});
notg #(0, 0) NOT_261 (c3540_wire_765, c3540_wire_83_3);
and_n #(2, 0, 0) AND_220 (c3540_wire_766, {c3540_wire_83_4, c3540_wire_767});
nor_n #(2, 0, 0) NOR_46 (c3540_wire_507, {c3540_wire_178_13, c3540_wire_150_17});
or_n #(2, 0, 0) OR_147 (c3540_wire_768, {c3540_wire_149_8, c3540_wire_151_10});
and_n #(3, 0, 0) AND_221 (c3540_wire_764, {c3540_wire_768, c3540_wire_506, c3540_wire_496});
or_n #(2, 0, 0) OR_148 (c3540_wire_84, {c3540_wire_769, c3540_wire_529});
notg #(0, 0) NOT_262 (c3540_wire_770, c3540_wire_84_2);
and_n #(2, 0, 0) AND_222 (c3540_wire_771, {c3540_wire_84_3, c3540_wire_772});
nor_n #(2, 0, 0) NOR_47 (c3540_wire_540, {c3540_wire_178_14, c3540_wire_150_18});
or_n #(2, 0, 0) OR_149 (c3540_wire_773, {c3540_wire_149_9, c3540_wire_151_11});
and_n #(3, 0, 0) AND_223 (c3540_wire_769, {c3540_wire_773, c3540_wire_539, c3540_wire_528});
nor_n #(2, 0, 0) NOR_48 (c3540_wire_774, {c3540_wire_112_1, c3540_wire_139});
or_n #(2, 0, 0) OR_150 (c3540_wire_775, {c3540_wire_136, c3540_wire_774});
notg #(0, 0) NOT_263 (c3540_wire_776, c3540_wire_694_0);
notg #(0, 0) NOT_264 (c3540_wire_777, c3540_wire_694_1);
notg #(0, 0) NOT_265 (c3540_wire_778, c3540_wire_715_0);
notg #(0, 0) NOT_266 (c3540_wire_779, c3540_wire_715_1);
notg #(0, 0) NOT_267 (c3540_wire_780, c3540_wire_733_0);
notg #(0, 0) NOT_268 (c3540_wire_781, c3540_wire_733_1);
or_n #(2, 0, 0) OR_151 (c3540_wire_782, {c3540_wire_733_2, c3540_wire_783});
or_n #(2, 0, 0) OR_152 (c3540_wire_784, {c3540_wire_738_0, c3540_wire_785_0});
and_n #(2, 0, 0) AND_224 (c3540_wire_159, {c3540_wire_150_19, c3540_wire_33_24});
bufg #(0, 0) BUF_18 (c3540_wire_149, G25_net_0);
or_n #(2, 0, 0) OR_153 (c3540_wire_740, {c3540_wire_786, c3540_wire_697});
notg #(0, 0) NOT_269 (c3540_wire_787, c3540_wire_740_2);
nor_n #(2, 0, 0) NOR_49 (c3540_wire_355, {c3540_wire_178_15, c3540_wire_150_20});
or_n #(2, 0, 0) OR_154 (c3540_wire_788, {c3540_wire_149_10, c3540_wire_151_12});
and_n #(3, 0, 0) AND_225 (c3540_wire_786, {c3540_wire_788, c3540_wire_696, c3540_wire_353});
or_n #(2, 0, 0) OR_155 (c3540_wire_85, {c3540_wire_789, c3540_wire_718});
notg #(0, 0) NOT_270 (c3540_wire_790, c3540_wire_85_2);
and_n #(2, 0, 0) AND_226 (c3540_wire_791, {c3540_wire_85_3, c3540_wire_792});
notg #(0, 0) NOT_271 (c3540_wire_793, c3540_wire_85_4);
or_n #(2, 0, 0) OR_156 (c3540_wire_794, {c3540_wire_85_5, c3540_wire_737});
nor_n #(2, 0, 0) NOR_50 (c3540_wire_474, {c3540_wire_178_16, c3540_wire_150_21});
or_n #(2, 0, 0) OR_157 (c3540_wire_795, {c3540_wire_149_11, c3540_wire_151_13});
and_n #(3, 0, 0) AND_227 (c3540_wire_789, {c3540_wire_795, c3540_wire_717, c3540_wire_472});
and_n #(2, 0, 0) AND_228 (c3540_wire_796, {c3540_wire_741_1, c3540_wire_797});
and_n #(4, 0, 0) AND_229 (c3540_wire_798, {c3540_wire_741_2, c3540_wire_799_0, c3540_wire_800_0, c3540_wire_732_1});
and_n #(2, 0, 0) AND_230 (c3540_wire_158, {c3540_wire_149_12, c3540_wire_33_25});
bufg #(0, 0) BUF_19 (c3540_wire_151, G26_net_0);
nand_n #(2, 0, 0) NAND_4 (c3540_wire_801, {c3540_wire_403_1, c3540_wire_742_3});
and_n #(2, 0, 0) AND_231 (c3540_wire_802, {c3540_wire_776, c3540_wire_803});
or_n #(2, 0, 0) OR_158 (c3540_wire_804, {c3540_wire_802, c3540_wire_745});
and_n #(2, 0, 0) AND_232 (c3540_wire_805, {c3540_wire_804, c3540_wire_729});
and_n #(2, 0, 0) AND_233 (c3540_wire_806, {c3540_wire_730, c3540_wire_801});
or_n #(2, 0, 0) OR_159 (c3540_wire_803, {c3540_wire_787, c3540_wire_806});
and_n #(2, 0, 0) AND_234 (c3540_wire_807, {c3540_wire_808, c3540_wire_734});
notg #(0, 0) NOT_272 (c3540_wire_797, c3540_wire_807_0);
nand_n #(2, 0, 0) NAND_5 (c3540_wire_809, {c3540_wire_525_2, c3540_wire_83_5});
or_n #(2, 0, 0) OR_160 (c3540_wire_810, {c3540_wire_793, c3540_wire_811});
and_n #(2, 0, 0) AND_235 (c3540_wire_812, {c3540_wire_810, c3540_wire_778});
or_n #(2, 0, 0) OR_161 (c3540_wire_808, {c3540_wire_812, c3540_wire_762});
and_n #(2, 0, 0) AND_236 (c3540_wire_811, {c3540_wire_735, c3540_wire_809});
notg #(0, 0) NOT_273 (c3540_wire_813, c3540_wire_805_0);
notg #(0, 0) NOT_274 (c3540_wire_814, c3540_wire_805_1);
nor_n #(2, 0, 0) NOR_51 (c3540_wire_815, {c3540_wire_807_1, c3540_wire_40_15});
notg #(0, 0) NOT_275 (c3540_wire_816, c3540_wire_815_0);
notg #(0, 0) NOT_276 (c3540_wire_817, c3540_wire_815_1);
notg #(0, 0) NOT_277 (c3540_wire_818, c3540_wire_815_2);
or_n #(2, 0, 0) OR_162 (c3540_wire_819, {c3540_wire_815_3, c3540_wire_820});
and_n #(2, 0, 0) AND_237 (c3540_wire_821, {c3540_wire_815_4, c3540_wire_588});
notg #(0, 0) NOT_278 (c3540_wire_822, c3540_wire_815_5);
or_n #(2, 0, 0) OR_163 (c3540_wire_823, {c3540_wire_815_6, c3540_wire_824_0});
xor_n #(2, 0, 0) XOR_8 (c3540_wire_825, {c3540_wire_815_7, c3540_wire_824_1});
notg #(0, 0) NOT_279 (c3540_wire_826, c3540_wire_827_0);
or_n #(2, 0, 0) OR_164 (c3540_wire_827, {c3540_wire_828, c3540_wire_81});
notg #(0, 0) NOT_280 (c3540_wire_829, c3540_wire_827_1);
notg #(0, 0) NOT_281 (c3540_wire_830, c3540_wire_827_2);
and_n #(2, 0, 0) AND_238 (c3540_wire_831, {c3540_wire_827_3, c3540_wire_832_0});
notg #(0, 0) NOT_282 (c3540_wire_833, c3540_wire_827_4);
or_n #(2, 0, 0) OR_165 (c3540_wire_834, {c3540_wire_453, c3540_wire_835});
and_n #(2, 0, 0) AND_239 (c3540_wire_828, {c3540_wire_834, c3540_wire_80});
nor_n #(5, 0, 0) NOR_52 (c3540_wire_835, {c3540_wire_454_4, c3540_wire_450_4, c3540_wire_455_4, c3540_wire_456_4, c3540_wire_150_22});
bufg #(0, 0) BUF_20 (c3540_wire_41, G27_net_0);
xor_n #(2, 0, 0) XOR_9 (c3540_wire_836, {c3540_wire_596_0, c3540_wire_837_0});
and_n #(2, 0, 0) AND_240 (c3540_wire_838, {c3540_wire_596_1, c3540_wire_60_32});
and_n #(2, 0, 0) AND_241 (c3540_wire_839, {c3540_wire_799_1, c3540_wire_780});
and_n #(2, 0, 0) AND_242 (c3540_wire_840, {c3540_wire_799_2, c3540_wire_732_2});
and_n #(2, 0, 0) AND_243 (c3540_wire_841, {c3540_wire_799_3, c3540_wire_800_1});
and_n #(2, 0, 0) AND_244 (c3540_wire_842, {c3540_wire_799_4, c3540_wire_732_3});
and_n #(2, 0, 0) AND_245 (c3540_wire_843, {c3540_wire_799_5, c3540_wire_732_4});
or_n #(2, 0, 0) OR_166 (c3540_wire_799, {c3540_wire_844, c3540_wire_749});
and_n #(2, 0, 0) AND_246 (c3540_wire_845, {c3540_wire_799_6, c3540_wire_60_33});
and_n #(2, 0, 0) AND_247 (c3540_wire_846, {c3540_wire_799_7, c3540_wire_830});
and_n #(2, 0, 0) AND_248 (c3540_wire_847, {c3540_wire_799_8, c3540_wire_848});
nand_n #(2, 0, 0) NAND_6 (c3540_wire_750, {c3540_wire_40_16, c3540_wire_73_4});
and_n #(2, 0, 0) AND_249 (c3540_wire_844, {c3540_wire_72, c3540_wire_748});
and_n #(2, 0, 0) AND_250 (c3540_wire_849, {c3540_wire_800_2, c3540_wire_826});
and_n #(2, 0, 0) AND_251 (c3540_wire_850, {c3540_wire_800_3, c3540_wire_817});
or_n #(2, 0, 0) OR_167 (c3540_wire_800, {c3540_wire_851, c3540_wire_754});
and_n #(2, 0, 0) AND_252 (c3540_wire_852, {c3540_wire_800_4, c3540_wire_60_34});
and_n #(2, 0, 0) AND_253 (c3540_wire_853, {c3540_wire_800_5, c3540_wire_832_1});
and_n #(2, 0, 0) AND_254 (c3540_wire_783, {c3540_wire_800_6, c3540_wire_818});
notg #(0, 0) NOT_283 (c3540_wire_820, c3540_wire_800_7);
and_n #(2, 0, 0) AND_255 (c3540_wire_854, {c3540_wire_800_8, c3540_wire_832_2});
nand_n #(2, 0, 0) NAND_7 (c3540_wire_755, {c3540_wire_40_17, c3540_wire_75_4});
and_n #(2, 0, 0) AND_256 (c3540_wire_851, {c3540_wire_74, c3540_wire_753});
or_n #(2, 0, 0) OR_168 (c3540_wire_855, {c3540_wire_856, c3540_wire_760});
and_n #(2, 0, 0) AND_257 (c3540_wire_857, {c3540_wire_855_0, c3540_wire_858});
notg #(0, 0) NOT_284 (c3540_wire_859, c3540_wire_855_1);
nand_n #(2, 0, 0) NAND_8 (c3540_wire_761, {c3540_wire_40_18, c3540_wire_69_4});
and_n #(2, 0, 0) AND_258 (c3540_wire_856, {c3540_wire_68, c3540_wire_759});
or_n #(2, 0, 0) OR_169 (c3540_wire_785, {c3540_wire_860, c3540_wire_766});
notg #(0, 0) NOT_285 (c3540_wire_861, c3540_wire_785_1);
notg #(0, 0) NOT_286 (c3540_wire_862, c3540_wire_785_2);
notg #(0, 0) NOT_287 (c3540_wire_863, c3540_wire_785_3);
nand_n #(2, 0, 0) NAND_9 (c3540_wire_767, {c3540_wire_40_19, c3540_wire_79_4});
and_n #(2, 0, 0) AND_259 (c3540_wire_860, {c3540_wire_78, c3540_wire_765});
or_n #(2, 0, 0) OR_170 (c3540_wire_864, {c3540_wire_865, c3540_wire_771});
and_n #(2, 0, 0) AND_260 (c3540_wire_866, {c3540_wire_864_0, c3540_wire_832_3});
and_n #(2, 0, 0) AND_261 (c3540_wire_867, {c3540_wire_864_1, c3540_wire_832_4});
and_n #(2, 0, 0) AND_262 (c3540_wire_868, {c3540_wire_864_2, c3540_wire_862});
notg #(0, 0) NOT_288 (c3540_wire_869, c3540_wire_864_3);
or_n #(2, 0, 0) OR_171 (c3540_wire_870, {c3540_wire_864_4, c3540_wire_871});
and_n #(2, 0, 0) AND_263 (c3540_wire_872, {c3540_wire_864_5, c3540_wire_832_5});
notg #(0, 0) NOT_289 (c3540_wire_873, c3540_wire_864_6);
nand_n #(2, 0, 0) NAND_10 (c3540_wire_772, {c3540_wire_40_20, c3540_wire_71_4});
and_n #(2, 0, 0) AND_264 (c3540_wire_865, {c3540_wire_70, c3540_wire_770});
or_n #(3, 0, 0) OR_172 (c3540_wire_874, {c3540_wire_170, c3540_wire_875, c3540_wire_876});
notg #(0, 0) NOT_290 (c3540_wire_877, c3540_wire_874);
notg #(0, 0) NOT_291 (c3540_wire_171, c3540_wire_18_9);
and_n #(2, 0, 0) AND_265 (c3540_wire_878, {c3540_wire_615, c3540_wire_60_35});
or_n #(2, 0, 0) OR_173 (c3540_wire_879, {c3540_wire_878, c3540_wire_880});
nor_n #(2, 0, 0) NOR_53 (c3540_wire_880, {c3540_wire_640, c3540_wire_60_36});
nor_n #(2, 0, 0) NOR_54 (c3540_wire_881, {c3540_wire_38_4, c3540_wire_18_10});
or_n #(2, 0, 0) OR_174 (c3540_wire_882, {c3540_wire_881, c3540_wire_883});
and_n #(2, 0, 0) AND_266 (c3540_wire_875, {c3540_wire_838, c3540_wire_884});
and_n #(2, 0, 0) AND_267 (c3540_wire_883, {c3540_wire_879, c3540_wire_38_5});
and_n #(2, 0, 0) AND_268 (c3540_wire_876, {c3540_wire_882, c3540_wire_169});
notg #(0, 0) NOT_292 (c3540_wire_884, c3540_wire_32_5);
and_n #(2, 0, 0) AND_269 (c3540_wire_885, {c3540_wire_732_5, c3540_wire_60_37});
and_n #(2, 0, 0) AND_270 (c3540_wire_886, {c3540_wire_732_6, c3540_wire_887});
or_n #(3, 0, 0) OR_175 (c3540_wire_888, {c3540_wire_889, c3540_wire_890, c3540_wire_167});
notg #(0, 0) NOT_293 (c3540_wire_891, c3540_wire_888);
notg #(0, 0) NOT_294 (c3540_wire_168, c3540_wire_121_14);
nor_n #(2, 0, 0) NOR_55 (c3540_wire_892, {c3540_wire_623, c3540_wire_60_38});
or_n #(2, 0, 0) OR_176 (c3540_wire_893, {c3540_wire_892, c3540_wire_894});
and_n #(2, 0, 0) AND_271 (c3540_wire_889, {c3540_wire_845, c3540_wire_895});
and_n #(2, 0, 0) AND_272 (c3540_wire_890, {c3540_wire_893, c3540_wire_166});
and_n #(2, 0, 0) AND_273 (c3540_wire_894, {c3540_wire_667, c3540_wire_60_39});
notg #(0, 0) NOT_295 (c3540_wire_895, c3540_wire_32_6);
or_n #(3, 0, 0) OR_177 (c3540_wire_896, {c3540_wire_897, c3540_wire_898, c3540_wire_173});
notg #(0, 0) NOT_296 (c3540_wire_899, c3540_wire_896);
nor_n #(2, 0, 0) NOR_56 (c3540_wire_900, {c3540_wire_630, c3540_wire_60_40});
or_n #(2, 0, 0) OR_178 (c3540_wire_901, {c3540_wire_900, c3540_wire_902});
and_n #(2, 0, 0) AND_274 (c3540_wire_897, {c3540_wire_852, c3540_wire_903});
and_n #(2, 0, 0) AND_275 (c3540_wire_898, {c3540_wire_901, c3540_wire_172});
and_n #(2, 0, 0) AND_276 (c3540_wire_902, {c3540_wire_680, c3540_wire_60_41});
notg #(0, 0) NOT_297 (c3540_wire_903, c3540_wire_32_7);
or_n #(2, 0, 0) OR_179 (c3540_wire_904, {c3540_wire_905, c3540_wire_791});
and_n #(2, 0, 0) AND_277 (c3540_wire_906, {c3540_wire_904_0, c3540_wire_907});
notg #(0, 0) NOT_298 (c3540_wire_908, c3540_wire_904_1);
nand_n #(2, 0, 0) NAND_11 (c3540_wire_792, {c3540_wire_40_21, c3540_wire_77_4});
and_n #(2, 0, 0) AND_278 (c3540_wire_905, {c3540_wire_76, c3540_wire_790});
or_n #(2, 0, 0) OR_180 (c3540_wire_909, {c3540_wire_736, c3540_wire_910});
and_n #(2, 0, 0) AND_279 (c3540_wire_911, {c3540_wire_909_0, c3540_wire_832_6});
and_n #(2, 0, 0) AND_280 (c3540_wire_912, {c3540_wire_909_1, c3540_wire_913_0});
and_n #(2, 0, 0) AND_281 (c3540_wire_914, {c3540_wire_909_2, c3540_wire_913_1});
nor_n #(2, 0, 0) NOR_57 (c3540_wire_910, {c3540_wire_785_4, c3540_wire_738_1});
notg #(0, 0) NOT_299 (c3540_wire_915, c3540_wire_41_5);
bufg #(0, 0) BUF_21 (c3540_wire_345, G28_net_0);
xor_n #(2, 0, 0) XOR_10 (c3540_wire_916, {c3540_wire_917_0, c3540_wire_837_1});
or_n #(2, 0, 0) OR_181 (c3540_wire_917, {c3540_wire_814, c3540_wire_918});
and_n #(2, 0, 0) AND_282 (c3540_wire_919, {c3540_wire_917_1, c3540_wire_832_7});
nor_n #(2, 0, 0) NOR_58 (c3540_wire_918, {c3540_wire_815_8, c3540_wire_741_3});
notg #(0, 0) NOT_300 (c3540_wire_920, c3540_wire_839);
and_n #(2, 0, 0) AND_283 (c3540_wire_921, {c3540_wire_841, c3540_wire_816});
notg #(0, 0) NOT_301 (c3540_wire_922, c3540_wire_921);
nor_n #(3, 0, 0) NOR_59 (c3540_wire_923, {c3540_wire_785_5, c3540_wire_904_2, c3540_wire_738_2});
notg #(0, 0) NOT_302 (c3540_wire_924, c3540_wire_923);
and_n #(2, 0, 0) AND_284 (c3540_wire_925, {c3540_wire_739, c3540_wire_86});
notg #(0, 0) NOT_303 (c3540_wire_926, c3540_wire_925);
or_n #(3, 0, 0) OR_182 (c3540_wire_927, {c3540_wire_928, c3540_wire_929, c3540_wire_175});
notg #(0, 0) NOT_304 (c3540_wire_930, c3540_wire_927);
notg #(0, 0) NOT_305 (c3540_wire_176, c3540_wire_120_10);
nor_n #(2, 0, 0) NOR_60 (c3540_wire_931, {c3540_wire_616, c3540_wire_60_42});
or_n #(2, 0, 0) OR_183 (c3540_wire_932, {c3540_wire_931, c3540_wire_933});
and_n #(2, 0, 0) AND_285 (c3540_wire_928, {c3540_wire_885, c3540_wire_934});
and_n #(2, 0, 0) AND_286 (c3540_wire_929, {c3540_wire_932, c3540_wire_174});
and_n #(2, 0, 0) AND_287 (c3540_wire_933, {c3540_wire_658, c3540_wire_60_43});
notg #(0, 0) NOT_306 (c3540_wire_934, c3540_wire_32_8);
and_n #(2, 0, 0) AND_288 (c3540_wire_935, {c3540_wire_853, c3540_wire_829});
and_n #(2, 0, 0) AND_289 (c3540_wire_936, {c3540_wire_935_0, c3540_wire_782_0});
and_n #(2, 0, 0) AND_290 (c3540_wire_937, {c3540_wire_935_1, c3540_wire_782_1});
and_n #(2, 0, 0) AND_291 (c3540_wire_938, {c3540_wire_866, c3540_wire_939});
xor_n #(2, 0, 0) XOR_11 (c3540_wire_858, {c3540_wire_938_0, c3540_wire_940_0});
xor_n #(2, 0, 0) XOR_12 (c3540_wire_941, {c3540_wire_938_1, c3540_wire_940_1});
nor_n #(2, 0, 0) NOR_61 (c3540_wire_939, {c3540_wire_785_6, c3540_wire_904_3});
and_n #(3, 0, 0) AND_292 (c3540_wire_942, {c3540_wire_922, c3540_wire_920, c3540_wire_87});
and_n #(2, 0, 0) AND_293 (c3540_wire_92, {c3540_wire_779, c3540_wire_794});
and_n #(2, 0, 0) AND_294 (c3540_wire_940, {c3540_wire_924, c3540_wire_91});
bufg #(0, 0) BUF_22 (c3540_wire_333, G29_net_0);
and_n #(2, 0, 0) AND_295 (c3540_wire_943, {c3540_wire_854, c3540_wire_846});
and_n #(2, 0, 0) AND_296 (c3540_wire_944, {c3540_wire_943_0, c3540_wire_942_0});
and_n #(2, 0, 0) AND_297 (c3540_wire_945, {c3540_wire_943_1, c3540_wire_942_1});
and_n #(2, 0, 0) AND_298 (c3540_wire_946, {c3540_wire_840, c3540_wire_849});
and_n #(2, 0, 0) AND_299 (c3540_wire_947, {c3540_wire_946_0, c3540_wire_832_8});
and_n #(2, 0, 0) AND_300 (c3540_wire_948, {c3540_wire_731, c3540_wire_89});
notg #(0, 0) NOT_307 (c3540_wire_949, c3540_wire_948);
and_n #(2, 0, 0) AND_301 (c3540_wire_950, {c3540_wire_842, c3540_wire_781});
and_n #(2, 0, 0) AND_302 (c3540_wire_951, {c3540_wire_843, c3540_wire_850});
and_n #(2, 0, 0) AND_303 (c3540_wire_952, {c3540_wire_784, c3540_wire_926});
nor_n #(3, 0, 0) NOR_62 (c3540_wire_953, {c3540_wire_40_22, c3540_wire_743_3, c3540_wire_807_2});
notg #(0, 0) NOT_308 (c3540_wire_954, c3540_wire_953);
and_n #(2, 0, 0) AND_304 (c3540_wire_913, {c3540_wire_867, c3540_wire_861});
or_n #(2, 0, 0) OR_184 (c3540_wire_955, {c3540_wire_48, c3540_wire_777});
and_n #(3, 0, 0) AND_305 (c3540_wire_837, {c3540_wire_949, c3540_wire_955, c3540_wire_956});
nor_n #(2, 0, 0) NOR_63 (c3540_wire_956, {c3540_wire_950, c3540_wire_951});
and_n #(2, 0, 0) AND_306 (c3540_wire_957, {c3540_wire_911, c3540_wire_868});
and_n #(2, 0, 0) AND_307 (c3540_wire_958, {c3540_wire_954, c3540_wire_819});
notg #(0, 0) NOT_309 (c3540_wire_959, c3540_wire_952_0);
and_n #(2, 0, 0) AND_308 (c3540_wire_960, {c3540_wire_952_1, c3540_wire_870});
notg #(0, 0) NOT_310 (c3540_wire_961, c3540_wire_32_9);
or_n #(2, 0, 0) OR_185 (c3540_wire_584, {c3540_wire_32_10, c3540_wire_962});
and_n #(2, 0, 0) AND_309 (c3540_wire_963, {c3540_wire_32_11, c3540_wire_33_26});
notg #(0, 0) NOT_311 (c3540_wire_964, c3540_wire_32_12);
notg #(0, 0) NOT_312 (c3540_wire_965, c3540_wire_32_13);
notg #(0, 0) NOT_313 (c3540_wire_966, c3540_wire_32_14);
notg #(0, 0) NOT_314 (c3540_wire_967, c3540_wire_32_15);
and_n #(2, 0, 0) AND_310 (c3540_wire_595, {c3540_wire_32_16, c3540_wire_33_27});
notg #(0, 0) NOT_315 (c3540_wire_968, c3540_wire_32_17);
and_n #(4, 0, 0) AND_311 (c3540_wire_969, {c3540_wire_32_18, c3540_wire_212, c3540_wire_203, c3540_wire_970});
bufg #(0, 0) BUF_23 (c3540_wire_33, G3_net_0);
bufg #(0, 0) BUF_24 (c3540_wire_9, G30_net_0);
nor_n #(3, 0, 0) NOR_64 (c3540_wire_971, {c3540_wire_18_11, c3540_wire_35_6, c3540_wire_119_1});
or_n #(2, 0, 0) OR_186 (c3540_wire_972, {c3540_wire_821, c3540_wire_971});
and_n #(2, 0, 0) AND_312 (c3540_wire_973, {c3540_wire_919, c3540_wire_974});
xor_n #(2, 0, 0) XOR_13 (c3540_wire_975, {c3540_wire_973_0, c3540_wire_976_0});
notg #(0, 0) NOT_316 (c3540_wire_977, c3540_wire_973_1);
or_n #(2, 0, 0) OR_187 (c3540_wire_978, {c3540_wire_973_2, c3540_wire_976_1});
nor_n #(2, 0, 0) NOR_65 (c3540_wire_974, {c3540_wire_827_5, c3540_wire_741_4});
notg #(0, 0) NOT_317 (c3540_wire_979, c3540_wire_958_0);
and_n #(2, 0, 0) AND_313 (c3540_wire_980, {c3540_wire_958_1, c3540_wire_981});
or_n #(2, 0, 0) OR_188 (c3540_wire_982, {c3540_wire_983, c3540_wire_980});
notg #(0, 0) NOT_318 (c3540_wire_984, c3540_wire_982);
nand_n #(2, 0, 0) NAND_12 (c3540_wire_981, {c3540_wire_827_6, c3540_wire_832_9});
and_n #(2, 0, 0) AND_314 (c3540_wire_983, {c3540_wire_831, c3540_wire_979});
bufg #(0, 0) BUF_25 (c3540_wire_10, G31_net_0);
or_n #(2, 0, 0) OR_189 (c3540_wire_985, {c3540_wire_872, c3540_wire_986});
nor_n #(2, 0, 0) NOR_66 (c3540_wire_986, {c3540_wire_864_7, c3540_wire_832_10});
nor_n #(2, 0, 0) NOR_67 (c3540_wire_987, {c3540_wire_5_13, c3540_wire_155_11});
nor_n #(2, 0, 0) NOR_68 (c3540_wire_988, {c3540_wire_157_14, c3540_wire_120_11});
nor_n #(2, 0, 0) NOR_69 (c3540_wire_989, {c3540_wire_161_15, c3540_wire_18_12});
notg #(0, 0) NOT_319 (c3540_wire_990, c3540_wire_60_44);
and_n #(2, 0, 0) AND_315 (c3540_wire_991, {c3540_wire_990, c3540_wire_992});
and_n #(2, 0, 0) AND_316 (c3540_wire_993, {c3540_wire_281, c3540_wire_994_0});
and_n #(2, 0, 0) AND_317 (c3540_wire_995, {c3540_wire_269, c3540_wire_549_3});
and_n #(2, 0, 0) AND_318 (c3540_wire_996, {c3540_wire_295, c3540_wire_997_0});
or_n #(2, 0, 0) OR_190 (c3540_wire_998, {c3540_wire_685_1, c3540_wire_999});
and_n #(2, 0, 0) AND_319 (c3540_wire_1000, {c3540_wire_998, c3540_wire_241});
or_n #(2, 0, 0) OR_191 (c3540_wire_1001, {c3540_wire_483_6, c3540_wire_1002_0});
and_n #(2, 0, 0) AND_320 (c3540_wire_1003, {c3540_wire_1001, c3540_wire_260});
and_n #(3, 0, 0) AND_321 (c3540_wire_1004, {c3540_wire_873, c3540_wire_1005, c3540_wire_60_45});
nor_n #(2, 0, 0) NOR_70 (c3540_wire_1006, {c3540_wire_32_19, c3540_wire_1_22});
nor_n #(2, 0, 0) NOR_71 (c3540_wire_1007, {c3540_wire_33_28, c3540_wire_469_5});
nand_n #(2, 0, 0) NAND_13 (c3540_wire_1008, {c3540_wire_35_7, c3540_wire_1009_0});
and_n #(2, 0, 0) AND_322 (c3540_wire_1010, {c3540_wire_1008, c3540_wire_985});
and_n #(2, 0, 0) AND_323 (c3540_wire_1011, {c3540_wire_728, c3540_wire_240});
nand_n #(2, 0, 0) NAND_14 (c3540_wire_1012, {c3540_wire_123_14, c3540_wire_121_15});
and_n #(2, 0, 0) AND_324 (c3540_wire_1013, {c3540_wire_1012, c3540_wire_259});
or_n #(2, 0, 0) OR_192 (c3540_wire_1014, {c3540_wire_987, c3540_wire_988});
or_n #(2, 0, 0) OR_193 (c3540_wire_992, {c3540_wire_989, c3540_wire_1015});
or_n #(5, 0, 0) OR_194 (c3540_wire_1005, {c3540_wire_993, c3540_wire_995, c3540_wire_996, c3540_wire_1000, c3540_wire_1003});
and_n #(3, 0, 0) AND_325 (c3540_wire_1016, {c3540_wire_1006, c3540_wire_1017, c3540_wire_38_6});
and_n #(2, 0, 0) AND_326 (c3540_wire_1018, {c3540_wire_1007, c3540_wire_1016});
or_n #(3, 0, 0) OR_195 (c3540_wire_1015, {c3540_wire_1011, c3540_wire_1013, c3540_wire_1014});
or_n #(2, 0, 0) OR_196 (c3540_wire_1019, {c3540_wire_1010, c3540_wire_1018});
or_n #(2, 0, 0) OR_197 (c3540_wire_1017, {c3540_wire_1004, c3540_wire_991});
or_n #(2, 0, 0) OR_198 (c3540_wire_887, {c3540_wire_944, c3540_wire_1020});
nor_n #(2, 0, 0) NOR_72 (c3540_wire_1020, {c3540_wire_943_2, c3540_wire_942_2});
or_n #(2, 0, 0) OR_199 (c3540_wire_1021, {c3540_wire_945, c3540_wire_1022});
or_n #(2, 0, 0) OR_200 (c3540_wire_1023, {c3540_wire_886, c3540_wire_1024});
nor_n #(2, 0, 0) NOR_73 (c3540_wire_1024, {c3540_wire_1021, c3540_wire_732_7});
nor_n #(2, 0, 0) NOR_74 (c3540_wire_1022, {c3540_wire_943_3, c3540_wire_942_3});
or_n #(2, 0, 0) OR_201 (c3540_wire_907, {c3540_wire_912, c3540_wire_1025});
nor_n #(2, 0, 0) NOR_75 (c3540_wire_1025, {c3540_wire_909_3, c3540_wire_913_2});
or_n #(2, 0, 0) OR_202 (c3540_wire_1026, {c3540_wire_914, c3540_wire_1027});
or_n #(2, 0, 0) OR_203 (c3540_wire_1028, {c3540_wire_906, c3540_wire_1029});
nor_n #(2, 0, 0) NOR_76 (c3540_wire_1029, {c3540_wire_1026, c3540_wire_904_4});
nor_n #(2, 0, 0) NOR_77 (c3540_wire_1027, {c3540_wire_909_4, c3540_wire_913_3});
and_n #(3, 0, 0) AND_327 (c3540_wire_1030, {c3540_wire_833, c3540_wire_1031, c3540_wire_832_11});
and_n #(2, 0, 0) AND_328 (c3540_wire_1032, {c3540_wire_1030_0, c3540_wire_916_0});
or_n #(2, 0, 0) OR_204 (c3540_wire_1031, {c3540_wire_798, c3540_wire_1033});
nor_n #(2, 0, 0) NOR_78 (c3540_wire_1033, {c3540_wire_741_5, c3540_wire_946_1});
or_n #(2, 0, 0) OR_205 (c3540_wire_824, {c3540_wire_1034, c3540_wire_960});
notg #(0, 0) NOT_320 (c3540_wire_871, c3540_wire_832_12);
and_n #(3, 0, 0) AND_329 (c3540_wire_1034, {c3540_wire_959, c3540_wire_869, c3540_wire_832_13});
notg #(0, 0) NOT_321 (c3540_wire_1035, c3540_wire_836_0);
and_n #(2, 0, 0) AND_330 (c3540_wire_1036, {c3540_wire_836_1, c3540_wire_1037});
and_n #(2, 0, 0) AND_331 (c3540_wire_1038, {c3540_wire_1023_0, c3540_wire_978});
and_n #(2, 0, 0) AND_332 (c3540_wire_1039, {c3540_wire_1028_0, c3540_wire_823});
or_n #(2, 0, 0) OR_206 (c3540_wire_1040, {c3540_wire_857, c3540_wire_1041});
notg #(0, 0) NOT_322 (c3540_wire_1042, c3540_wire_1040);
nor_n #(2, 0, 0) NOR_79 (c3540_wire_1041, {c3540_wire_855_2, c3540_wire_941});
nand_n #(2, 0, 0) NAND_15 (c3540_wire_1043, {c3540_wire_35_8, c3540_wire_1009_1});
and_n #(2, 0, 0) AND_333 (c3540_wire_1044, {c3540_wire_984, c3540_wire_1043});
or_n #(2, 0, 0) OR_207 (c3540_wire_1045, {c3540_wire_1044, c3540_wire_1046});
and_n #(6, 0, 0) AND_334 (c3540_wire_1046, {c3540_wire_964, c3540_wire_589, c3540_wire_899, c3540_wire_1047, c3540_wire_1048, c3540_wire_38_7});
notg #(0, 0) NOT_323 (c3540_wire_1047, c3540_wire_33_29);
notg #(0, 0) NOT_324 (c3540_wire_1048, c3540_wire_1049_0);
and_n #(2, 0, 0) AND_335 (c3540_wire_22, {c3540_wire_10_5, c3540_wire_1050});
bufg #(0, 0) BUF_26 (c3540_wire_401, G32_net_0);
or_n #(2, 0, 0) OR_208 (c3540_wire_976, {c3540_wire_847, c3540_wire_1051});
or_n #(2, 0, 0) OR_209 (c3540_wire_848, {c3540_wire_936, c3540_wire_1052});
or_n #(2, 0, 0) OR_210 (c3540_wire_1053, {c3540_wire_937, c3540_wire_1054});
nor_n #(2, 0, 0) NOR_80 (c3540_wire_1051, {c3540_wire_1053, c3540_wire_799_9});
nor_n #(2, 0, 0) NOR_81 (c3540_wire_1052, {c3540_wire_935_2, c3540_wire_782_2});
nor_n #(2, 0, 0) NOR_82 (c3540_wire_1054, {c3540_wire_935_3, c3540_wire_782_3});
or_n #(2, 0, 0) OR_211 (c3540_wire_1055, {c3540_wire_1032, c3540_wire_1056});
and_n #(2, 0, 0) AND_336 (c3540_wire_1057, {c3540_wire_968, c3540_wire_1058});
notg #(0, 0) NOT_325 (c3540_wire_970, c3540_wire_33_30);
and_n #(2, 0, 0) AND_337 (c3540_wire_1059, {c3540_wire_593, c3540_wire_1060});
and_n #(2, 0, 0) AND_338 (c3540_wire_1061, {c3540_wire_594, c3540_wire_1055});
nor_n #(2, 0, 0) NOR_83 (c3540_wire_1056, {c3540_wire_1030_1, c3540_wire_916_1});
and_n #(2, 0, 0) AND_339 (c3540_wire_1062, {c3540_wire_1063, c3540_wire_18_13});
or_n #(2, 0, 0) OR_212 (c3540_wire_1058, {c3540_wire_1062, c3540_wire_1064});
and_n #(2, 0, 0) AND_340 (c3540_wire_1065, {c3540_wire_1066, c3540_wire_1067});
or_n #(2, 0, 0) OR_213 (c3540_wire_1068, {c3540_wire_1065, c3540_wire_1069});
nor_n #(2, 0, 0) NOR_84 (c3540_wire_1069, {c3540_wire_120_12, c3540_wire_121_16});
or_n #(2, 0, 0) OR_214 (c3540_wire_1060, {c3540_wire_969, c3540_wire_1057});
and_n #(2, 0, 0) AND_341 (c3540_wire_1064, {c3540_wire_1068, c3540_wire_63});
or_n #(2, 0, 0) OR_215 (c3540_wire_1070, {c3540_wire_1061, c3540_wire_1059});
notg #(0, 0) NOT_326 (c3540_wire_1063, c3540_wire_121_17);
and_n #(2, 0, 0) AND_342 (c3540_wire_1066, {c3540_wire_120_13, c3540_wire_121_18});
notg #(0, 0) NOT_327 (c3540_wire_1067, c3540_wire_18_14);
or_n #(2, 0, 0) OR_216 (c3540_wire_1071, {c3540_wire_1072, c3540_wire_1036});
notg #(0, 0) NOT_328 (c3540_wire_1073, c3540_wire_1071);
nand_n #(2, 0, 0) NAND_16 (c3540_wire_1037, {c3540_wire_946_2, c3540_wire_832_14});
and_n #(2, 0, 0) AND_343 (c3540_wire_1072, {c3540_wire_947, c3540_wire_1035});
nor_n #(2, 0, 0) NOR_85 (c3540_wire_1074, {c3540_wire_824_2, c3540_wire_1028_1});
and_n #(2, 0, 0) AND_344 (c3540_wire_1075, {c3540_wire_253, c3540_wire_725});
nor_n #(2, 0, 0) NOR_86 (c3540_wire_1076, {c3540_wire_155_12, c3540_wire_120_14});
notg #(0, 0) NOT_329 (c3540_wire_1077, c3540_wire_60_46);
and_n #(2, 0, 0) AND_345 (c3540_wire_1078, {c3540_wire_1077, c3540_wire_1079});
and_n #(2, 0, 0) AND_346 (c3540_wire_1080, {c3540_wire_290, c3540_wire_685_2});
and_n #(2, 0, 0) AND_347 (c3540_wire_1081, {c3540_wire_277, c3540_wire_549_4});
or_n #(2, 0, 0) OR_217 (c3540_wire_1082, {c3540_wire_483_7, c3540_wire_1002_1});
and_n #(2, 0, 0) AND_348 (c3540_wire_1083, {c3540_wire_1082, c3540_wire_235});
or_n #(2, 0, 0) OR_218 (c3540_wire_1084, {c3540_wire_135, c3540_wire_516_4});
or_n #(2, 0, 0) OR_219 (c3540_wire_1085, {c3540_wire_822, c3540_wire_1074});
and_n #(2, 0, 0) AND_349 (c3540_wire_1086, {c3540_wire_254, c3540_wire_1084});
nor_n #(2, 0, 0) NOR_87 (c3540_wire_1087, {c3540_wire_181_13, c3540_wire_155_13});
and_n #(3, 0, 0) AND_350 (c3540_wire_1088, {c3540_wire_859, c3540_wire_1089, c3540_wire_60_47});
nor_n #(2, 0, 0) NOR_88 (c3540_wire_1090, {c3540_wire_32_20, c3540_wire_1_23});
nor_n #(2, 0, 0) NOR_89 (c3540_wire_1091, {c3540_wire_33_31, c3540_wire_469_6});
or_n #(2, 0, 0) OR_220 (c3540_wire_1092, {c3540_wire_690, c3540_wire_608});
and_n #(2, 0, 0) AND_351 (c3540_wire_1093, {c3540_wire_143, c3540_wire_1085});
and_n #(2, 0, 0) AND_352 (c3540_wire_1094, {c3540_wire_580, c3540_wire_234});
or_n #(3, 0, 0) OR_221 (c3540_wire_1079, {c3540_wire_1076, c3540_wire_1092, c3540_wire_1095});
or_n #(2, 0, 0) OR_222 (c3540_wire_1096, {c3540_wire_1080, c3540_wire_1081});
or_n #(2, 0, 0) OR_223 (c3540_wire_1097, {c3540_wire_1083, c3540_wire_1086});
or_n #(3, 0, 0) OR_224 (c3540_wire_1089, {c3540_wire_1087, c3540_wire_1096, c3540_wire_1097});
and_n #(3, 0, 0) AND_353 (c3540_wire_1098, {c3540_wire_1090, c3540_wire_1099, c3540_wire_38_8});
notg #(0, 0) NOT_330 (c3540_wire_1100, c3540_wire_1009_2);
or_n #(2, 0, 0) OR_225 (c3540_wire_1101, {c3540_wire_1100, c3540_wire_1093});
and_n #(2, 0, 0) AND_354 (c3540_wire_1102, {c3540_wire_1091, c3540_wire_1098});
or_n #(2, 0, 0) OR_226 (c3540_wire_1095, {c3540_wire_1094, c3540_wire_1075});
and_n #(2, 0, 0) AND_355 (c3540_wire_1103, {c3540_wire_1042, c3540_wire_1101});
or_n #(2, 0, 0) OR_227 (c3540_wire_1104, {c3540_wire_1103, c3540_wire_1102});
or_n #(2, 0, 0) OR_228 (c3540_wire_1099, {c3540_wire_1078, c3540_wire_1088});
notg #(0, 0) NOT_331 (c3540_wire_581, c3540_wire_18_15);
and_n #(2, 0, 0) AND_356 (c3540_wire_1105, {c3540_wire_825, c3540_wire_145});
nor_n #(2, 0, 0) NOR_90 (c3540_wire_1106, {c3540_wire_157_15, c3540_wire_18_16});
notg #(0, 0) NOT_332 (c3540_wire_1107, c3540_wire_60_48);
and_n #(2, 0, 0) AND_357 (c3540_wire_1108, {c3540_wire_1107, c3540_wire_1109});
and_n #(2, 0, 0) AND_358 (c3540_wire_1110, {c3540_wire_280, c3540_wire_1002_2});
and_n #(2, 0, 0) AND_359 (c3540_wire_1111, {c3540_wire_268, c3540_wire_516_5});
and_n #(2, 0, 0) AND_360 (c3540_wire_1112, {c3540_wire_294, c3540_wire_994_1});
or_n #(2, 0, 0) OR_229 (c3540_wire_1113, {c3540_wire_549_5, c3540_wire_997_1});
and_n #(2, 0, 0) AND_361 (c3540_wire_1114, {c3540_wire_1113, c3540_wire_239});
or_n #(2, 0, 0) OR_230 (c3540_wire_1115, {c3540_wire_213, c3540_wire_685_3});
and_n #(2, 0, 0) AND_362 (c3540_wire_1116, {c3540_wire_258, c3540_wire_1115});
and_n #(3, 0, 0) AND_363 (c3540_wire_1117, {c3540_wire_863, c3540_wire_1118, c3540_wire_60_49});
nor_n #(2, 0, 0) NOR_91 (c3540_wire_1119, {c3540_wire_32_21, c3540_wire_1_24});
nor_n #(2, 0, 0) NOR_92 (c3540_wire_1120, {c3540_wire_33_32, c3540_wire_469_7});
nor_n #(2, 0, 0) NOR_93 (c3540_wire_1121, {c3540_wire_824_3, c3540_wire_1009_3});
or_n #(3, 0, 0) OR_231 (c3540_wire_1122, {c3540_wire_1105, c3540_wire_1121, c3540_wire_1123});
or_n #(5, 0, 0) OR_232 (c3540_wire_1109, {c3540_wire_727, c3540_wire_1124, c3540_wire_1106, c3540_wire_1125, c3540_wire_1126});
and_n #(2, 0, 0) AND_364 (c3540_wire_1125, {c3540_wire_692, c3540_wire_238});
notg #(0, 0) NOT_333 (c3540_wire_693, c3540_wire_121_19);
nand_n #(2, 0, 0) NAND_17 (c3540_wire_1127, {c3540_wire_99_15, c3540_wire_120_15});
and_n #(2, 0, 0) AND_365 (c3540_wire_1126, {c3540_wire_1127, c3540_wire_257});
nor_n #(2, 0, 0) NOR_94 (c3540_wire_1124, {c3540_wire_2_16, c3540_wire_155_14});
or_n #(4, 0, 0) OR_233 (c3540_wire_1128, {c3540_wire_1110, c3540_wire_1111, c3540_wire_1112, c3540_wire_1114});
and_n #(3, 0, 0) AND_366 (c3540_wire_1129, {c3540_wire_1119, c3540_wire_1130, c3540_wire_38_9});
and_n #(2, 0, 0) AND_367 (c3540_wire_1123, {c3540_wire_1120, c3540_wire_1129});
or_n #(2, 0, 0) OR_234 (c3540_wire_1118, {c3540_wire_1128, c3540_wire_1116});
or_n #(2, 0, 0) OR_235 (c3540_wire_1130, {c3540_wire_1108, c3540_wire_1117});
nor_n #(3, 0, 0) NOR_95 (c3540_wire_1131, {c3540_wire_824_4, c3540_wire_815_9, c3540_wire_1028_2});
nand_n #(2, 0, 0) NAND_18 (c3540_wire_1132, {c3540_wire_18_17, c3540_wire_5_14});
and_n #(2, 0, 0) AND_368 (c3540_wire_1133, {c3540_wire_255, c3540_wire_1132});
nor_n #(2, 0, 0) NOR_96 (c3540_wire_1134, {c3540_wire_155_15, c3540_wire_121_20});
notg #(0, 0) NOT_334 (c3540_wire_1135, c3540_wire_60_50);
and_n #(2, 0, 0) AND_369 (c3540_wire_1136, {c3540_wire_1135, c3540_wire_1137});
and_n #(2, 0, 0) AND_370 (c3540_wire_1138, {c3540_wire_279, c3540_wire_685_4});
and_n #(2, 0, 0) AND_371 (c3540_wire_1139, {c3540_wire_267, c3540_wire_483_8});
and_n #(2, 0, 0) AND_372 (c3540_wire_1140, {c3540_wire_292, c3540_wire_1002_3});
or_n #(2, 0, 0) OR_236 (c3540_wire_1141, {c3540_wire_516_6, c3540_wire_994_2});
and_n #(2, 0, 0) AND_373 (c3540_wire_1142, {c3540_wire_1141, c3540_wire_237});
or_n #(2, 0, 0) OR_237 (c3540_wire_1143, {c3540_wire_191, c3540_wire_549_6});
and_n #(2, 0, 0) AND_374 (c3540_wire_1144, {c3540_wire_256, c3540_wire_1143});
and_n #(3, 0, 0) AND_375 (c3540_wire_1145, {c3540_wire_908, c3540_wire_1146, c3540_wire_60_51});
nor_n #(2, 0, 0) NOR_97 (c3540_wire_1147, {c3540_wire_32_22, c3540_wire_1_25});
nor_n #(2, 0, 0) NOR_98 (c3540_wire_1148, {c3540_wire_33_33, c3540_wire_469_8});
nor_n #(2, 0, 0) NOR_99 (c3540_wire_1149, {c3540_wire_1028_3, c3540_wire_1009_4});
or_n #(2, 0, 0) OR_238 (c3540_wire_1150, {c3540_wire_1039, c3540_wire_1131});
or_n #(2, 0, 0) OR_239 (c3540_wire_1151, {c3540_wire_726, c3540_wire_691});
and_n #(2, 0, 0) AND_376 (c3540_wire_1152, {c3540_wire_609, c3540_wire_236});
or_n #(3, 0, 0) OR_240 (c3540_wire_1137, {c3540_wire_1134, c3540_wire_1151, c3540_wire_1153});
or_n #(4, 0, 0) OR_241 (c3540_wire_1154, {c3540_wire_1138, c3540_wire_1139, c3540_wire_1140, c3540_wire_1142});
and_n #(2, 0, 0) AND_377 (c3540_wire_1155, {c3540_wire_144, c3540_wire_1150});
and_n #(3, 0, 0) AND_378 (c3540_wire_1156, {c3540_wire_1147, c3540_wire_1157, c3540_wire_38_10});
and_n #(2, 0, 0) AND_379 (c3540_wire_1158, {c3540_wire_1148, c3540_wire_1156});
or_n #(3, 0, 0) OR_242 (c3540_wire_1159, {c3540_wire_1149, c3540_wire_1155, c3540_wire_1158});
or_n #(2, 0, 0) OR_243 (c3540_wire_1153, {c3540_wire_1152, c3540_wire_1133});
or_n #(2, 0, 0) OR_244 (c3540_wire_1146, {c3540_wire_1154, c3540_wire_1144});
or_n #(2, 0, 0) OR_245 (c3540_wire_1157, {c3540_wire_1145, c3540_wire_1136});
notg #(0, 0) NOT_335 (c3540_wire_610, c3540_wire_120_16);
and_n #(2, 0, 0) AND_380 (c3540_wire_23, {c3540_wire_401_7, c3540_wire_1160});
bufg #(0, 0) BUF_27 (c3540_wire_430, G33_net_0);
nor_n #(3, 0, 0) NOR_100 (c3540_wire_1161, {c3540_wire_1023_1, c3540_wire_973_3, c3540_wire_976_2});
nor_n #(2, 0, 0) NOR_101 (c3540_wire_1162, {c3540_wire_1023_2, c3540_wire_1009_5});
or_n #(2, 0, 0) OR_246 (c3540_wire_1163, {c3540_wire_1038, c3540_wire_1161});
and_n #(6, 0, 0) AND_381 (c3540_wire_1164, {c3540_wire_967, c3540_wire_592, c3540_wire_930, c3540_wire_1165, c3540_wire_1166, c3540_wire_38_11});
or_n #(3, 0, 0) OR_247 (c3540_wire_1167, {c3540_wire_1164, c3540_wire_1162, c3540_wire_1168});
and_n #(2, 0, 0) AND_382 (c3540_wire_1168, {c3540_wire_1163, c3540_wire_142});
notg #(0, 0) NOT_336 (c3540_wire_1165, c3540_wire_33_34);
notg #(0, 0) NOT_337 (c3540_wire_1166, c3540_wire_1049_1);
and_n #(2, 0, 0) AND_383 (c3540_wire_1169, {c3540_wire_975, c3540_wire_140});
and_n #(6, 0, 0) AND_384 (c3540_wire_1170, {c3540_wire_965, c3540_wire_590, c3540_wire_891, c3540_wire_1171, c3540_wire_1172, c3540_wire_38_12});
or_n #(3, 0, 0) OR_248 (c3540_wire_1173, {c3540_wire_1170, c3540_wire_1174, c3540_wire_1169});
nor_n #(2, 0, 0) NOR_102 (c3540_wire_1174, {c3540_wire_976_3, c3540_wire_1009_6});
notg #(0, 0) NOT_338 (c3540_wire_1171, c3540_wire_33_35);
notg #(0, 0) NOT_339 (c3540_wire_1172, c3540_wire_1049_2);
nor_n #(2, 0, 0) NOR_103 (c3540_wire_1175, {c3540_wire_1023_3, c3540_wire_976_4});
notg #(0, 0) NOT_340 (c3540_wire_1176, c3540_wire_1049_3);
and_n #(6, 0, 0) AND_385 (c3540_wire_1177, {c3540_wire_1176, c3540_wire_966, c3540_wire_591, c3540_wire_877, c3540_wire_1178, c3540_wire_38_13});
or_n #(2, 0, 0) OR_249 (c3540_wire_1179, {c3540_wire_1175, c3540_wire_977});
or_n #(2, 0, 0) OR_250 (c3540_wire_1180, {c3540_wire_1177, c3540_wire_1181});
and_n #(2, 0, 0) AND_386 (c3540_wire_1182, {c3540_wire_1179, c3540_wire_141});
or_n #(2, 0, 0) OR_251 (c3540_wire_1183, {c3540_wire_1182, c3540_wire_1184});
and_n #(2, 0, 0) AND_387 (c3540_wire_1181, {c3540_wire_1183, c3540_wire_1073});
notg #(0, 0) NOT_341 (c3540_wire_1184, c3540_wire_1009_7);
notg #(0, 0) NOT_342 (c3540_wire_1178, c3540_wire_33_36);
and_n #(2, 0, 0) AND_388 (c3540_wire_1185, {c3540_wire_1019_0, c3540_wire_1122_0});
or_n #(2, 0, 0) OR_252 (c3540_wire_1186, {c3540_wire_1185, c3540_wire_1187});
nor_n #(2, 0, 0) NOR_104 (c3540_wire_1187, {c3540_wire_1122_1, c3540_wire_1019_1});
notg #(0, 0) NOT_343 (c3540_wire_1188, c3540_wire_1189);
nor_n #(8, 0, 0) NOR_105 (c3540_wire_1189, {c3540_wire_1019_2, c3540_wire_1122_2, c3540_wire_1159_0, c3540_wire_1104_0, c3540_wire_1045_0, c3540_wire_1173_0, c3540_wire_1167_0, c3540_wire_1180_0});
and_n #(2, 0, 0) AND_389 (c3540_wire_1190, {c3540_wire_1186_0, c3540_wire_1191});
and_n #(2, 0, 0) AND_390 (c3540_wire_24, {c3540_wire_430_7, c3540_wire_49});
bufg #(0, 0) BUF_28 (c3540_wire_28, G34_net_0);
and_n #(2, 0, 0) AND_391 (c3540_wire_1192, {c3540_wire_1167_1, c3540_wire_1180_1});
or_n #(2, 0, 0) OR_253 (c3540_wire_1193, {c3540_wire_1192, c3540_wire_1194});
nor_n #(2, 0, 0) NOR_106 (c3540_wire_1194, {c3540_wire_1180_2, c3540_wire_1167_2});
xor_n #(2, 0, 0) XOR_14 (c3540_wire_1195, {c3540_wire_1045_1, c3540_wire_1173_1});
xor_n #(2, 0, 0) XOR_15 (c3540_wire_195, {c3540_wire_1195_0, c3540_wire_1196_0});
xor_n #(2, 0, 0) XOR_16 (c3540_wire_1197, {c3540_wire_1195_1, c3540_wire_1196_1});
and_n #(2, 0, 0) AND_392 (c3540_wire_1198, {c3540_wire_1195_2, c3540_wire_1199});
xor_n #(2, 0, 0) XOR_17 (c3540_wire_1199, {c3540_wire_1193_0, c3540_wire_1200_0});
xor_n #(2, 0, 0) XOR_18 (c3540_wire_1201, {c3540_wire_1193_1, c3540_wire_1200_1});
and_n #(2, 0, 0) AND_393 (c3540_wire_1196, {c3540_wire_1202, c3540_wire_95});
xor_n #(2, 0, 0) XOR_19 (c3540_wire_1202, {c3540_wire_1167_3, c3540_wire_1180_3});
xor_n #(2, 0, 0) XOR_20 (c3540_wire_1203, {c3540_wire_1200_2, c3540_wire_1204});
or_n #(2, 0, 0) OR_254 (c3540_wire_1200, {c3540_wire_1190, c3540_wire_1205});
and_n #(2, 0, 0) AND_394 (c3540_wire_1206, {c3540_wire_1104_1, c3540_wire_1159_1});
or_n #(2, 0, 0) OR_255 (c3540_wire_1191, {c3540_wire_1206, c3540_wire_1207});
or_n #(2, 0, 0) OR_256 (c3540_wire_1208, {c3540_wire_1209, c3540_wire_1210});
nor_n #(2, 0, 0) NOR_107 (c3540_wire_1205, {c3540_wire_1208, c3540_wire_1186_1});
nor_n #(2, 0, 0) NOR_108 (c3540_wire_1207, {c3540_wire_1104_2, c3540_wire_1159_2});
and_n #(2, 0, 0) AND_395 (c3540_wire_1209, {c3540_wire_1104_3, c3540_wire_1159_3});
nor_n #(2, 0, 0) NOR_109 (c3540_wire_1210, {c3540_wire_1104_4, c3540_wire_1159_4});
or_n #(2, 0, 0) OR_257 (c3540_wire_1204, {c3540_wire_194, c3540_wire_1211});
nor_n #(2, 0, 0) NOR_110 (c3540_wire_1211, {c3540_wire_192_1, c3540_wire_1197});
bufg #(0, 0) BUF_29 (c3540_wire_111, G35_net_0);
nor_n #(2, 0, 0) NOR_111 (c3540_wire_1212, {c3540_wire_1195_3, c3540_wire_1201});
or_n #(2, 0, 0) OR_258 (c3540_wire_1213, {c3540_wire_1198, c3540_wire_1212});
bufg #(0, 0) BUF_30 (G3519_net_0, c3540_wire_1214);
and_n #(2, 0, 0) AND_396 (c3540_wire_1214, {c3540_wire_309_1, c3540_wire_50});
bufg #(0, 0) BUF_31 (G3520_net_0, c3540_wire_6);
bufg #(0, 0) BUF_32 (G3521_net_0, c3540_wire_558);
bufg #(0, 0) BUF_33 (G3522_net_0, c3540_wire_775);
bufg #(0, 0) BUF_34 (G3523_net_0, c3540_wire_1215);
or_n #(2, 0, 0) OR_259 (c3540_wire_219, {c3540_wire_220, c3540_wire_1216});
or_n #(2, 0, 0) OR_260 (c3540_wire_1217, {c3540_wire_222, c3540_wire_1218});
or_n #(2, 0, 0) OR_261 (c3540_wire_1215, {c3540_wire_218, c3540_wire_1219});
nor_n #(2, 0, 0) NOR_112 (c3540_wire_1219, {c3540_wire_1217, c3540_wire_198_1});
nor_n #(2, 0, 0) NOR_113 (c3540_wire_1216, {c3540_wire_200_2, c3540_wire_221_2});
nor_n #(2, 0, 0) NOR_114 (c3540_wire_1218, {c3540_wire_200_3, c3540_wire_221_3});
bufg #(0, 0) BUF_35 (G3524_net_0, c3540_wire_758);
bufg #(0, 0) BUF_36 (G3525_net_0, c3540_wire_1220);
or_n #(2, 0, 0) OR_262 (c3540_wire_1220, {c3540_wire_813, c3540_wire_796});
bufg #(0, 0) BUF_37 (G3526_net_0, c3540_wire_957);
bufg #(0, 0) BUF_38 (G3527_net_0, c3540_wire_972);
bufg #(0, 0) BUF_39 (G3528_net_0, c3540_wire_1019_3);
bufg #(0, 0) BUF_40 (G3529_net_0, c3540_wire_1045_2);
bufg #(0, 0) BUF_41 (G3530_net_0, c3540_wire_1070);
bufg #(0, 0) BUF_42 (G3531_net_0, c3540_wire_1104_5);
bufg #(0, 0) BUF_43 (G3532_net_0, c3540_wire_1122_3);
bufg #(0, 0) BUF_44 (G3533_net_0, c3540_wire_1159_5);
bufg #(0, 0) BUF_45 (G3534_net_0, c3540_wire_1167_4);
notg #(0, 0) NOT_344 (c3540_wire_1221, c3540_wire_1167_5);
bufg #(0, 0) BUF_46 (G3535_net_0, c3540_wire_1180_4);
notg #(0, 0) NOT_345 (c3540_wire_1222, c3540_wire_1180_5);
bufg #(0, 0) BUF_47 (G3536_net_0, c3540_wire_1173_2);
bufg #(0, 0) BUF_48 (G3537_net_0, c3540_wire_1188);
bufg #(0, 0) BUF_49 (G3538_net_0, c3540_wire_1223);
nor_n #(6, 0, 0) NOR_115 (c3540_wire_97, {c3540_wire_1045_3, c3540_wire_1019_4, c3540_wire_1104_6, c3540_wire_1159_6, c3540_wire_1122_4, c3540_wire_1173_3});
and_n #(3, 0, 0) AND_397 (c3540_wire_1224, {c3540_wire_96, c3540_wire_1222, c3540_wire_1221});
or_n #(2, 0, 0) OR_263 (c3540_wire_1223, {c3540_wire_1224, c3540_wire_915});
bufg #(0, 0) BUF_50 (G3539_net_0, c3540_wire_1203);
bufg #(0, 0) BUF_51 (G3540_net_0, c3540_wire_1213);
and_n #(2, 0, 0) AND_398 (c3540_wire_25, {c3540_wire_111_6, c3540_wire_124});
bufg #(0, 0) BUF_52 (c3540_wire_115, G36_net_0);
and_n #(2, 0, 0) AND_399 (c3540_wire_26, {c3540_wire_115_5, c3540_wire_179});
bufg #(0, 0) BUF_53 (c3540_wire_116, G37_net_0);
and_n #(2, 0, 0) AND_400 (c3540_wire_27, {c3540_wire_116_3, c3540_wire_204});
bufg #(0, 0) BUF_54 (c3540_wire_340, G38_net_0);
bufg #(0, 0) BUF_55 (c3540_wire_483, G39_net_0);
and_n #(2, 0, 0) AND_401 (c3540_wire_326, {c3540_wire_33_37, c3540_wire_582});
notg #(0, 0) NOT_346 (c3540_wire_1225, c3540_wire_33_38);
and_n #(2, 0, 0) AND_402 (c3540_wire_962, {c3540_wire_33_39, c3540_wire_60_52});
bufg #(0, 0) BUF_56 (c3540_wire_60, G4_net_0);
bufg #(0, 0) BUF_57 (c3540_wire_516, G40_net_0);
bufg #(0, 0) BUF_58 (c3540_wire_549, G41_net_0);
bufg #(0, 0) BUF_59 (c3540_wire_685, G42_net_0);
bufg #(0, 0) BUF_60 (c3540_wire_1002, G43_net_0);
bufg #(0, 0) BUF_61 (c3540_wire_994, G44_net_0);
bufg #(0, 0) BUF_62 (c3540_wire_997, G45_net_0);
bufg #(0, 0) BUF_63 (c3540_wire_999, G46_net_0);
bufg #(0, 0) BUF_64 (c3540_wire_832, G47_net_0);
bufg #(0, 0) BUF_65 (c3540_wire_42, G48_net_0);
bufg #(0, 0) BUF_66 (c3540_wire_344, G49_net_0);
and_n #(2, 0, 0) AND_403 (c3540_wire_449, {c3540_wire_60_53, c3540_wire_583});
bufg #(0, 0) BUF_67 (c3540_wire_38, G5_net_0);
bufg #(0, 0) BUF_68 (c3540_wire_193, G50_net_0);
or_n #(2, 0, 0) OR_264 (c3540_wire_1226, {c3540_wire_38_14, c3540_wire_469_9});
bufg #(0, 0) BUF_69 (c3540_wire_469, G6_net_0);
and_n #(3, 0, 0) AND_404 (c3540_wire_1049, {c3540_wire_469_10, c3540_wire_1225, c3540_wire_961});
bufg #(0, 0) BUF_70 (c3540_wire_18, G7_net_0);
nor_n #(3, 0, 0) NOR_116 (c3540_wire_309, {c3540_wire_120_17, c3540_wire_18_18, c3540_wire_121_21});
notg #(0, 0) NOT_347 (c3540_wire_1050, c3540_wire_120_18);
notg #(0, 0) NOT_348 (c3540_wire_1160, c3540_wire_121_22);
and_n #(2, 0, 0) AND_405 (c3540_wire_341, {c3540_wire_1226, c3540_wire_585});
nor_n #(3, 0, 0) NOR_117 (c3540_wire_492, {c3540_wire_469_11, c3540_wire_1_26, c3540_wire_38_15});
nor_n #(3, 0, 0) NOR_118 (c3540_wire_441, {c3540_wire_99_16, c3540_wire_5_15, c3540_wire_123_15});
bufg #(0, 0) BUF_71 (c3540_wire_120, G8_net_0);
and_n #(2, 0, 0) AND_406 (c3540_wire_318, {c3540_wire_963, c3540_wire_586});
bufg #(0, 0) BUF_72 (c3540_wire_121, G9_net_0);
nor_n #(2, 0, 0) NOR_119 (c3540_wire_1009, {c3540_wire_1_27, c3540_wire_1049_4});
and_n #(2, 0, 0) AND_407 (c3540_wire_346, {c3540_wire_587, c3540_wire_1227});
nand_n #(2, 0, 0) NAND_19 (c3540_wire_1227, {c3540_wire_60_54, c3540_wire_38_16});

endmodule
