module Fictitious_DSP(Input, Output);

	input [15:0] Input;
	output [3:0] Output;

	// Fictitious DSP

endmodule