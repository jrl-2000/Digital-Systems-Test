
//Verilog file of module c1908


`timescale 1 ns / 1ns

module c1908_net(G1,
G10,
G11,
G12,
G13,
G14,
G15,
G16,
G17,
G18,
G1884,
G1885,
G1886,
G1887,
G1888,
G1889,
G1890,
G1891,
G1892,
G1893,
G1894,
G1895,
G1896,
G1897,
G1898,
G1899,
G19,
G1900,
G1901,
G1902,
G1903,
G1904,
G1905,
G1906,
G1907,
G1908,
G2,
G20,
G21,
G22,
G23,
G24,
G25,
G26,
G27,
G28,
G29,
G3,
G30,
G31,
G32,
G33,
G4,
G5,
G6,
G7,
G8,
G9);
input G1;
input G2;
input G3;
input G4;
input G5;
input G6;
input G7;
input G8;
input G9;
input G10;
input G11;
input G12;
input G13;
input G14;
input G15;
input G16;
input G17;
input G18;
input G19;
input G20;
input G21;
input G22;
input G23;
input G24;
input G25;
input G26;
input G27;
input G28;
input G29;
input G30;
input G31;
input G32;
input G33;

output G1884;
output G1885;
output G1886;
output G1887;
output G1888;
output G1889;
output G1890;
output G1891;
output G1892;
output G1893;
output G1894;
output G1895;
output G1896;
output G1897;
output G1898;
output G1899;
output G1900;
output G1901;
output G1902;
output G1903;
output G1904;
output G1905;
output G1906;
output G1907;
output G1908;

wire
c1908_wire_1,
c1908_wire_2,
c1908_wire_3,
c1908_wire_4,
c1908_wire_5,
c1908_wire_6,
c1908_wire_7,
c1908_wire_8,
c1908_wire_9,
c1908_wire_10,
c1908_wire_11,
c1908_wire_12,
c1908_wire_13,
c1908_wire_14,
c1908_wire_15,
c1908_wire_16,
c1908_wire_17,
c1908_wire_18,
c1908_wire_19,
c1908_wire_20,
c1908_wire_21,
c1908_wire_22,
c1908_wire_23,
c1908_wire_24,
c1908_wire_25,
c1908_wire_26,
c1908_wire_27,
c1908_wire_28,
c1908_wire_29,
c1908_wire_30,
c1908_wire_31,
c1908_wire_32,
c1908_wire_33,
c1908_wire_34,
c1908_wire_35,
c1908_wire_36,
c1908_wire_37,
c1908_wire_38,
c1908_wire_39,
c1908_wire_40,
c1908_wire_41,
c1908_wire_42,
c1908_wire_43,
c1908_wire_44,
c1908_wire_45,
c1908_wire_46,
c1908_wire_47,
c1908_wire_48,
c1908_wire_49,
c1908_wire_50,
c1908_wire_51,
c1908_wire_52,
c1908_wire_53,
c1908_wire_54,
c1908_wire_55,
c1908_wire_56,
c1908_wire_57,
c1908_wire_58,
c1908_wire_59,
c1908_wire_60,
c1908_wire_61,
c1908_wire_62,
c1908_wire_63,
c1908_wire_64,
c1908_wire_65,
c1908_wire_66,
c1908_wire_67,
c1908_wire_68,
c1908_wire_69,
c1908_wire_70,
c1908_wire_71,
c1908_wire_72,
c1908_wire_73,
c1908_wire_74,
c1908_wire_75,
c1908_wire_76,
c1908_wire_77,
c1908_wire_78,
c1908_wire_79,
c1908_wire_80,
c1908_wire_81,
c1908_wire_82,
c1908_wire_83,
c1908_wire_84,
c1908_wire_85,
c1908_wire_86,
c1908_wire_87,
c1908_wire_88,
c1908_wire_89,
c1908_wire_90,
c1908_wire_91,
c1908_wire_92,
c1908_wire_93,
c1908_wire_94,
c1908_wire_95,
c1908_wire_96,
c1908_wire_97,
c1908_wire_98,
c1908_wire_99,
c1908_wire_100,
c1908_wire_101,
c1908_wire_102,
c1908_wire_103,
c1908_wire_104,
c1908_wire_105,
c1908_wire_106,
c1908_wire_107,
c1908_wire_108,
c1908_wire_109,
c1908_wire_110,
c1908_wire_111,
c1908_wire_112,
c1908_wire_113,
c1908_wire_114,
c1908_wire_115,
c1908_wire_116,
c1908_wire_117,
c1908_wire_118,
c1908_wire_119,
c1908_wire_120,
c1908_wire_121,
c1908_wire_122,
c1908_wire_123,
c1908_wire_124,
c1908_wire_125,
c1908_wire_126,
c1908_wire_127,
c1908_wire_128,
c1908_wire_129,
c1908_wire_130,
c1908_wire_131,
c1908_wire_132,
c1908_wire_133,
c1908_wire_134,
c1908_wire_135,
c1908_wire_136,
c1908_wire_137,
c1908_wire_138,
c1908_wire_139,
c1908_wire_140,
c1908_wire_141,
c1908_wire_142,
c1908_wire_143,
c1908_wire_144,
c1908_wire_145,
c1908_wire_146,
c1908_wire_147,
c1908_wire_148,
c1908_wire_149,
c1908_wire_150,
c1908_wire_151,
c1908_wire_152,
c1908_wire_153,
c1908_wire_154,
c1908_wire_155,
c1908_wire_156,
c1908_wire_157,
c1908_wire_158,
c1908_wire_159,
c1908_wire_160,
c1908_wire_161,
c1908_wire_162,
c1908_wire_163,
c1908_wire_164,
c1908_wire_165,
c1908_wire_166,
c1908_wire_167,
c1908_wire_168,
c1908_wire_169,
c1908_wire_170,
c1908_wire_171,
c1908_wire_172,
c1908_wire_173,
c1908_wire_174,
c1908_wire_175,
c1908_wire_176,
c1908_wire_177,
c1908_wire_178,
c1908_wire_179,
c1908_wire_180,
c1908_wire_181,
c1908_wire_182,
c1908_wire_183,
c1908_wire_184,
c1908_wire_185,
c1908_wire_186,
c1908_wire_187,
c1908_wire_188,
c1908_wire_189,
c1908_wire_190,
c1908_wire_191,
c1908_wire_192,
c1908_wire_193,
c1908_wire_194,
c1908_wire_195,
c1908_wire_196,
c1908_wire_197,
c1908_wire_198,
c1908_wire_199,
c1908_wire_200,
c1908_wire_201,
c1908_wire_202,
c1908_wire_203,
c1908_wire_204,
c1908_wire_205,
c1908_wire_206,
c1908_wire_207,
c1908_wire_208,
c1908_wire_209,
c1908_wire_210,
c1908_wire_211,
c1908_wire_212,
c1908_wire_213,
c1908_wire_214,
c1908_wire_215,
c1908_wire_216,
c1908_wire_217,
c1908_wire_218,
c1908_wire_219,
c1908_wire_220,
c1908_wire_221,
c1908_wire_222,
c1908_wire_223,
c1908_wire_224,
c1908_wire_225,
c1908_wire_226,
c1908_wire_227,
c1908_wire_228,
c1908_wire_229,
c1908_wire_230,
c1908_wire_231,
c1908_wire_232,
c1908_wire_233,
c1908_wire_234,
c1908_wire_235,
c1908_wire_236,
c1908_wire_237,
c1908_wire_238,
c1908_wire_239,
c1908_wire_240,
c1908_wire_241,
c1908_wire_242,
c1908_wire_243,
c1908_wire_244,
c1908_wire_245,
c1908_wire_246,
c1908_wire_247,
c1908_wire_248,
c1908_wire_249,
c1908_wire_250,
c1908_wire_251,
c1908_wire_252,
c1908_wire_253,
c1908_wire_254,
c1908_wire_255,
c1908_wire_256,
c1908_wire_257,
c1908_wire_258,
c1908_wire_259,
c1908_wire_260,
c1908_wire_261,
c1908_wire_262,
c1908_wire_263,
c1908_wire_264,
c1908_wire_265,
c1908_wire_266,
c1908_wire_267,
c1908_wire_268,
c1908_wire_269,
c1908_wire_270,
c1908_wire_271,
c1908_wire_272,
c1908_wire_273,
c1908_wire_274,
c1908_wire_275,
c1908_wire_276,
c1908_wire_277,
c1908_wire_278,
c1908_wire_279,
c1908_wire_280,
c1908_wire_281,
c1908_wire_282,
c1908_wire_283,
c1908_wire_284,
c1908_wire_285,
c1908_wire_286,
c1908_wire_287,
c1908_wire_288,
c1908_wire_289,
c1908_wire_290,
c1908_wire_291,
c1908_wire_292,
c1908_wire_293,
c1908_wire_294,
c1908_wire_295,
c1908_wire_296,
c1908_wire_297,
c1908_wire_298,
c1908_wire_299,
c1908_wire_300,
c1908_wire_301,
c1908_wire_302,
c1908_wire_303,
c1908_wire_304,
c1908_wire_305,
c1908_wire_306,
c1908_wire_307,
c1908_wire_308,
c1908_wire_309,
c1908_wire_310,
c1908_wire_311,
c1908_wire_312,
c1908_wire_313,
c1908_wire_314,
c1908_wire_315,
c1908_wire_316,
c1908_wire_317,
c1908_wire_318,
c1908_wire_319,
c1908_wire_320,
c1908_wire_321,
c1908_wire_322,
c1908_wire_323,
c1908_wire_324,
c1908_wire_325,
c1908_wire_326,
c1908_wire_327,
c1908_wire_328,
c1908_wire_329,
c1908_wire_330,
c1908_wire_331,
c1908_wire_332,
c1908_wire_333,
c1908_wire_334,
c1908_wire_335,
c1908_wire_336,
c1908_wire_337,
c1908_wire_338,
c1908_wire_339,
c1908_wire_340,
c1908_wire_341,
c1908_wire_342,
c1908_wire_343,
c1908_wire_344,
c1908_wire_345,
c1908_wire_346,
c1908_wire_347,
c1908_wire_348,
c1908_wire_349,
c1908_wire_350,
c1908_wire_351,
c1908_wire_352,
c1908_wire_353,
c1908_wire_354,
c1908_wire_355,
c1908_wire_356,
c1908_wire_357,
c1908_wire_358,
c1908_wire_359,
c1908_wire_360,
c1908_wire_361,
c1908_wire_362,
c1908_wire_363,
c1908_wire_364,
c1908_wire_365,
c1908_wire_366,
c1908_wire_367,
c1908_wire_368,
c1908_wire_369,
c1908_wire_370,
c1908_wire_371,
c1908_wire_372,
c1908_wire_373,
c1908_wire_374,
c1908_wire_375,
c1908_wire_376,
c1908_wire_377,
c1908_wire_378,
c1908_wire_379,
c1908_wire_380,
c1908_wire_381,
c1908_wire_382,
c1908_wire_383,
c1908_wire_384,
c1908_wire_385,
c1908_wire_386,
c1908_wire_387,
c1908_wire_388,
c1908_wire_389,
c1908_wire_390,
c1908_wire_391,
c1908_wire_392,
c1908_wire_393,
c1908_wire_394,
c1908_wire_395,
c1908_wire_396,
c1908_wire_397,
c1908_wire_398,
c1908_wire_399,
c1908_wire_400,
c1908_wire_401,
c1908_wire_402,
c1908_wire_403,
c1908_wire_404,
c1908_wire_405,
c1908_wire_406,
c1908_wire_407,
c1908_wire_408,
c1908_wire_409,
c1908_wire_410,
c1908_wire_411,
c1908_wire_412,
c1908_wire_413,
c1908_wire_414,
c1908_wire_415,
c1908_wire_416,
c1908_wire_417,
c1908_wire_418,
c1908_wire_419,
c1908_wire_420,
c1908_wire_421,
c1908_wire_422,
c1908_wire_423,
c1908_wire_424,
c1908_wire_425,
c1908_wire_426,
c1908_wire_427,
c1908_wire_428,
c1908_wire_429,
c1908_wire_430,
c1908_wire_431,
c1908_wire_432,
c1908_wire_433,
c1908_wire_434,
c1908_wire_1_0,
c1908_wire_1_1,
c1908_wire_1_2,
c1908_wire_1_3,
c1908_wire_1_4,
c1908_wire_2_0,
c1908_wire_2_1,
c1908_wire_2_2,
c1908_wire_2_3,
c1908_wire_2_4,
c1908_wire_2_5,
c1908_wire_2_6,
c1908_wire_2_7,
c1908_wire_4_0,
c1908_wire_4_1,
c1908_wire_4_2,
c1908_wire_4_3,
c1908_wire_14_0,
c1908_wire_14_1,
c1908_wire_5_0,
c1908_wire_5_1,
c1908_wire_5_2,
c1908_wire_5_3,
c1908_wire_5_4,
c1908_wire_17_0,
c1908_wire_17_1,
c1908_wire_17_2,
c1908_wire_17_3,
c1908_wire_34_0,
c1908_wire_34_1,
c1908_wire_34_2,
c1908_wire_34_3,
c1908_wire_45_0,
c1908_wire_45_1,
c1908_wire_45_2,
c1908_wire_45_3,
c1908_wire_60_0,
c1908_wire_60_1,
c1908_wire_60_2,
c1908_wire_60_3,
c1908_wire_31_0,
c1908_wire_31_1,
c1908_wire_31_2,
c1908_wire_31_3,
c1908_wire_31_4,
c1908_wire_31_5,
c1908_wire_82_0,
c1908_wire_82_1,
c1908_wire_82_2,
c1908_wire_93_0,
c1908_wire_93_1,
c1908_wire_93_2,
c1908_wire_29_0,
c1908_wire_29_1,
c1908_wire_29_2,
c1908_wire_29_3,
c1908_wire_29_4,
c1908_wire_29_5,
c1908_wire_35_0,
c1908_wire_35_1,
c1908_wire_35_2,
c1908_wire_35_3,
c1908_wire_35_4,
c1908_wire_35_5,
c1908_wire_35_6,
c1908_wire_115_0,
c1908_wire_115_1,
c1908_wire_115_2,
c1908_wire_49_0,
c1908_wire_49_1,
c1908_wire_49_2,
c1908_wire_49_3,
c1908_wire_121_0,
c1908_wire_121_1,
c1908_wire_121_2,
c1908_wire_121_3,
c1908_wire_135_0,
c1908_wire_135_1,
c1908_wire_125_0,
c1908_wire_125_1,
c1908_wire_125_2,
c1908_wire_125_3,
c1908_wire_125_4,
c1908_wire_140_0,
c1908_wire_140_1,
c1908_wire_140_2,
c1908_wire_30_0,
c1908_wire_30_1,
c1908_wire_30_2,
c1908_wire_30_3,
c1908_wire_30_4,
c1908_wire_30_5,
c1908_wire_151_0,
c1908_wire_151_1,
c1908_wire_151_2,
c1908_wire_151_3,
c1908_wire_151_4,
c1908_wire_151_5,
c1908_wire_151_6,
c1908_wire_151_7,
c1908_wire_151_8,
c1908_wire_151_9,
c1908_wire_155_0,
c1908_wire_155_1,
c1908_wire_155_2,
c1908_wire_155_3,
c1908_wire_155_4,
c1908_wire_155_5,
c1908_wire_155_6,
c1908_wire_155_7,
c1908_wire_155_8,
c1908_wire_155_9,
c1908_wire_185_0,
c1908_wire_185_1,
c1908_wire_156_0,
c1908_wire_156_1,
c1908_wire_156_2,
c1908_wire_156_3,
c1908_wire_156_4,
c1908_wire_156_5,
c1908_wire_156_6,
c1908_wire_156_7,
c1908_wire_156_8,
c1908_wire_156_9,
c1908_wire_200_0,
c1908_wire_200_1,
c1908_wire_200_2,
c1908_wire_200_3,
c1908_wire_211_0,
c1908_wire_211_1,
c1908_wire_211_2,
c1908_wire_211_3,
c1908_wire_211_4,
c1908_wire_67_0,
c1908_wire_67_1,
c1908_wire_67_2,
c1908_wire_67_3,
c1908_wire_67_4,
c1908_wire_67_5,
c1908_wire_67_6,
c1908_wire_157_0,
c1908_wire_157_1,
c1908_wire_157_2,
c1908_wire_157_3,
c1908_wire_157_4,
c1908_wire_157_5,
c1908_wire_157_6,
c1908_wire_157_7,
c1908_wire_157_8,
c1908_wire_157_9,
c1908_wire_167_0,
c1908_wire_167_1,
c1908_wire_167_2,
c1908_wire_167_3,
c1908_wire_167_4,
c1908_wire_167_5,
c1908_wire_167_6,
c1908_wire_233_0,
c1908_wire_233_1,
c1908_wire_233_2,
c1908_wire_233_3,
c1908_wire_233_4,
c1908_wire_233_5,
c1908_wire_56_0,
c1908_wire_56_1,
c1908_wire_21_0,
c1908_wire_21_1,
c1908_wire_21_2,
c1908_wire_21_3,
c1908_wire_21_4,
c1908_wire_21_5,
c1908_wire_21_6,
c1908_wire_21_7,
c1908_wire_241_0,
c1908_wire_241_1,
c1908_wire_241_2,
c1908_wire_241_3,
c1908_wire_241_4,
c1908_wire_22_0,
c1908_wire_22_1,
c1908_wire_22_2,
c1908_wire_22_3,
c1908_wire_22_4,
c1908_wire_22_5,
c1908_wire_161_0,
c1908_wire_161_1,
c1908_wire_161_2,
c1908_wire_258_0,
c1908_wire_258_1,
c1908_wire_258_2,
c1908_wire_258_3,
c1908_wire_258_4,
c1908_wire_258_5,
c1908_wire_258_6,
c1908_wire_258_7,
c1908_wire_258_8,
c1908_wire_258_9,
c1908_wire_70_0,
c1908_wire_70_1,
c1908_wire_70_2,
c1908_wire_70_3,
c1908_wire_70_4,
c1908_wire_70_5,
c1908_wire_70_6,
c1908_wire_218_0,
c1908_wire_218_1,
c1908_wire_218_2,
c1908_wire_218_3,
c1908_wire_218_4,
c1908_wire_218_5,
c1908_wire_218_6,
c1908_wire_277_0,
c1908_wire_277_1,
c1908_wire_277_2,
c1908_wire_277_3,
c1908_wire_277_4,
c1908_wire_277_5,
c1908_wire_277_6,
c1908_wire_277_7,
c1908_wire_277_8,
c1908_wire_277_9,
c1908_wire_287_0,
c1908_wire_287_1,
c1908_wire_287_2,
c1908_wire_101_0,
c1908_wire_101_1,
c1908_wire_101_2,
c1908_wire_101_3,
c1908_wire_101_4,
c1908_wire_101_5,
c1908_wire_101_6,
c1908_wire_101_7,
c1908_wire_101_8,
c1908_wire_290_0,
c1908_wire_290_1,
c1908_wire_290_2,
c1908_wire_290_3,
c1908_wire_291_0,
c1908_wire_291_1,
c1908_wire_291_2,
c1908_wire_291_3,
c1908_wire_291_4,
c1908_wire_291_5,
c1908_wire_235_0,
c1908_wire_235_1,
c1908_wire_235_2,
c1908_wire_235_3,
c1908_wire_235_4,
c1908_wire_302_0,
c1908_wire_302_1,
c1908_wire_302_2,
c1908_wire_302_3,
c1908_wire_137_0,
c1908_wire_137_1,
c1908_wire_203_0,
c1908_wire_203_1,
c1908_wire_318_0,
c1908_wire_318_1,
c1908_wire_318_2,
c1908_wire_318_3,
c1908_wire_252_0,
c1908_wire_252_1,
c1908_wire_197_0,
c1908_wire_197_1,
c1908_wire_197_2,
c1908_wire_197_3,
c1908_wire_197_4,
c1908_wire_79_0,
c1908_wire_79_1,
c1908_wire_143_0,
c1908_wire_143_1,
c1908_wire_143_2,
c1908_wire_143_3,
c1908_wire_143_4,
c1908_wire_11_0,
c1908_wire_11_1,
c1908_wire_11_2,
c1908_wire_11_3,
c1908_wire_11_4,
c1908_wire_11_5,
c1908_wire_408_0,
c1908_wire_408_1,
c1908_wire_169_0,
c1908_wire_169_1,
c1908_wire_169_2,
c1908_wire_169_3,
c1908_wire_169_4,
c1908_wire_169_5,
c1908_wire_169_6,
c1908_wire_213_0,
c1908_wire_213_1,
c1908_wire_85_0,
c1908_wire_85_1,
c1908_wire_85_2,
c1908_wire_52_0,
c1908_wire_52_1,
c1908_wire_52_2,
c1908_wire_52_3,
c1908_wire_52_4,
c1908_wire_52_5,
c1908_wire_193_0,
c1908_wire_193_1,
c1908_wire_193_2,
c1908_wire_193_3,
c1908_wire_193_4,
c1908_wire_193_5,
c1908_wire_193_6,
c1908_wire_300_0,
c1908_wire_300_1,
c1908_wire_300_2,
c1908_wire_300_3,
c1908_wire_300_4,
c1908_wire_413_0,
c1908_wire_413_1,
c1908_wire_413_2,
c1908_wire_231_0,
c1908_wire_231_1,
c1908_wire_231_2,
c1908_wire_216_0,
c1908_wire_216_1,
c1908_wire_216_2,
c1908_wire_183_0,
c1908_wire_183_1,
c1908_wire_183_2,
c1908_wire_172_0,
c1908_wire_172_1,
c1908_wire_172_2,
c1908_wire_150_0,
c1908_wire_150_1,
c1908_wire_150_2,
c1908_wire_12_0,
c1908_wire_12_1,
c1908_wire_12_2,
c1908_wire_12_3,
c1908_wire_12_4,
c1908_wire_12_5,
c1908_wire_387_0,
c1908_wire_387_1,
c1908_wire_387_2,
c1908_wire_96_0,
c1908_wire_96_1,
c1908_wire_96_2,
c1908_wire_96_3,
c1908_wire_96_4,
c1908_wire_96_5,
c1908_wire_96_6,
c1908_wire_96_7,
c1908_wire_96_8,
c1908_wire_96_9,
c1908_wire_96_10,
c1908_wire_96_11,
c1908_wire_96_12,
c1908_wire_96_13,
c1908_wire_96_14,
c1908_wire_96_15,
c1908_wire_96_16,
c1908_wire_96_17,
c1908_wire_96_18,
c1908_wire_96_19,
c1908_wire_96_20,
c1908_wire_361_0,
c1908_wire_361_1,
c1908_wire_361_2,
c1908_wire_365_0,
c1908_wire_365_1,
c1908_wire_365_2,
c1908_wire_365_3,
c1908_wire_365_4,
c1908_wire_365_5,
c1908_wire_54_0,
c1908_wire_54_1,
c1908_wire_54_2,
c1908_wire_54_3,
c1908_wire_54_4,
c1908_wire_54_5,
c1908_wire_54_6,
c1908_wire_54_7,
c1908_wire_54_8,
c1908_wire_54_9,
c1908_wire_54_10,
c1908_wire_54_11,
c1908_wire_54_12,
c1908_wire_54_13,
c1908_wire_54_14,
c1908_wire_54_15,
c1908_wire_54_16,
c1908_wire_54_17,
c1908_wire_54_18,
c1908_wire_237_0,
c1908_wire_237_1,
c1908_wire_237_2,
c1908_wire_237_3,
c1908_wire_239_0,
c1908_wire_239_1,
c1908_wire_239_2,
c1908_wire_239_3,
c1908_wire_239_4,
c1908_wire_239_5,
c1908_wire_239_6,
c1908_wire_303_0,
c1908_wire_303_1,
c1908_wire_303_2,
c1908_wire_303_3,
c1908_wire_43_0,
c1908_wire_43_1,
c1908_wire_43_2,
c1908_wire_43_3,
c1908_wire_43_4,
c1908_wire_43_5,
c1908_wire_163_0,
c1908_wire_163_1,
c1908_wire_163_2,
c1908_wire_163_3,
c1908_wire_163_4,
c1908_wire_41_0,
c1908_wire_41_1,
c1908_wire_41_2,
c1908_wire_41_3,
c1908_wire_41_4,
c1908_wire_41_5,
c1908_wire_42_0,
c1908_wire_42_1,
c1908_wire_42_2,
c1908_wire_42_3,
c1908_wire_42_4,
c1908_wire_42_5,
c1908_wire_36_0,
c1908_wire_36_1,
c1908_wire_106_0,
c1908_wire_106_1,
c1908_wire_106_2,
c1908_wire_106_3,
c1908_wire_106_4,
c1908_wire_111_0,
c1908_wire_111_1,
c1908_wire_265_0,
c1908_wire_265_1,
c1908_wire_265_2,
c1908_wire_268_0,
c1908_wire_268_1,
c1908_wire_268_2,
c1908_wire_279_0,
c1908_wire_279_1,
c1908_wire_279_2,
c1908_wire_279_3,
c1908_wire_279_4,
c1908_wire_279_5,
c1908_wire_279_6,
c1908_wire_279_7,
c1908_wire_15_0,
c1908_wire_15_1,
c1908_wire_15_2,
c1908_wire_15_3,
c1908_wire_15_4,
c1908_wire_15_5,
c1908_wire_15_6,
c1908_wire_112_0,
c1908_wire_112_1,
c1908_wire_87_0,
c1908_wire_87_1,
c1908_wire_87_2,
c1908_wire_87_3,
c1908_wire_88_0,
c1908_wire_88_1,
c1908_wire_88_2,
c1908_wire_88_3,
c1908_wire_76_0,
c1908_wire_76_1,
c1908_wire_77_0,
c1908_wire_77_1,
G1_net_0,
G2_net_0,
G3_net_0,
G4_net_0,
G5_net_0,
G6_net_0,
G7_net_0,
G8_net_0,
G9_net_0,
G10_net_0,
G11_net_0,
G12_net_0,
G13_net_0,
G14_net_0,
G15_net_0,
G16_net_0,
G17_net_0,
G18_net_0,
G19_net_0,
G20_net_0,
G21_net_0,
G22_net_0,
G23_net_0,
G24_net_0,
G25_net_0,
G26_net_0,
G27_net_0,
G28_net_0,
G29_net_0,
G30_net_0,
G31_net_0,
G32_net_0,
G33_net_0,
G1884_net_0,
G1885_net_0,
G1886_net_0,
G1887_net_0,
G1888_net_0,
G1889_net_0,
G1890_net_0,
G1891_net_0,
G1892_net_0,
G1893_net_0,
G1894_net_0,
G1895_net_0,
G1896_net_0,
G1897_net_0,
G1898_net_0,
G1899_net_0,
G1900_net_0,
G1901_net_0,
G1902_net_0,
G1903_net_0,
G1904_net_0,
G1905_net_0,
G1906_net_0,
G1907_net_0,
G1908_net_0;

pin #(33) pin_0 ({G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33}, {G1_net_0, G2_net_0, G3_net_0, G4_net_0, G5_net_0, G6_net_0, G7_net_0, G8_net_0, G9_net_0, G10_net_0, G11_net_0, G12_net_0, G13_net_0, G14_net_0, G15_net_0, G16_net_0, G17_net_0, G18_net_0, G19_net_0, G20_net_0, G21_net_0, G22_net_0, G23_net_0, G24_net_0, G25_net_0, G26_net_0, G27_net_0, G28_net_0, G29_net_0, G30_net_0, G31_net_0, G32_net_0, G33_net_0});

pout #(25) pout_0 ({G1884_net_0, G1885_net_0, G1886_net_0, G1887_net_0, G1888_net_0, G1889_net_0, G1890_net_0, G1891_net_0, G1892_net_0, G1893_net_0, G1894_net_0, G1895_net_0, G1896_net_0, G1897_net_0, G1898_net_0, G1899_net_0, G1900_net_0, G1901_net_0, G1902_net_0, G1903_net_0, G1904_net_0, G1905_net_0, G1906_net_0, G1907_net_0, G1908_net_0}, {G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893, G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903, G1904, G1905, G1906, G1907, G1908});

fanout_n #(5, 0, 0) FANOUT_1 (c1908_wire_1, {c1908_wire_1_0, c1908_wire_1_1, c1908_wire_1_2, c1908_wire_1_3, c1908_wire_1_4});
fanout_n #(8, 0, 0) FANOUT_2 (c1908_wire_2, {c1908_wire_2_0, c1908_wire_2_1, c1908_wire_2_2, c1908_wire_2_3, c1908_wire_2_4, c1908_wire_2_5, c1908_wire_2_6, c1908_wire_2_7});
fanout_n #(4, 0, 0) FANOUT_3 (c1908_wire_4, {c1908_wire_4_0, c1908_wire_4_1, c1908_wire_4_2, c1908_wire_4_3});
fanout_n #(2, 0, 0) FANOUT_4 (c1908_wire_14, {c1908_wire_14_0, c1908_wire_14_1});
fanout_n #(5, 0, 0) FANOUT_5 (c1908_wire_5, {c1908_wire_5_0, c1908_wire_5_1, c1908_wire_5_2, c1908_wire_5_3, c1908_wire_5_4});
fanout_n #(4, 0, 0) FANOUT_6 (c1908_wire_17, {c1908_wire_17_0, c1908_wire_17_1, c1908_wire_17_2, c1908_wire_17_3});
fanout_n #(4, 0, 0) FANOUT_7 (c1908_wire_34, {c1908_wire_34_0, c1908_wire_34_1, c1908_wire_34_2, c1908_wire_34_3});
fanout_n #(4, 0, 0) FANOUT_8 (c1908_wire_45, {c1908_wire_45_0, c1908_wire_45_1, c1908_wire_45_2, c1908_wire_45_3});
fanout_n #(4, 0, 0) FANOUT_9 (c1908_wire_60, {c1908_wire_60_0, c1908_wire_60_1, c1908_wire_60_2, c1908_wire_60_3});
fanout_n #(6, 0, 0) FANOUT_10 (c1908_wire_31, {c1908_wire_31_0, c1908_wire_31_1, c1908_wire_31_2, c1908_wire_31_3, c1908_wire_31_4, c1908_wire_31_5});
fanout_n #(3, 0, 0) FANOUT_11 (c1908_wire_82, {c1908_wire_82_0, c1908_wire_82_1, c1908_wire_82_2});
fanout_n #(3, 0, 0) FANOUT_12 (c1908_wire_93, {c1908_wire_93_0, c1908_wire_93_1, c1908_wire_93_2});
fanout_n #(6, 0, 0) FANOUT_13 (c1908_wire_29, {c1908_wire_29_0, c1908_wire_29_1, c1908_wire_29_2, c1908_wire_29_3, c1908_wire_29_4, c1908_wire_29_5});
fanout_n #(7, 0, 0) FANOUT_14 (c1908_wire_35, {c1908_wire_35_0, c1908_wire_35_1, c1908_wire_35_2, c1908_wire_35_3, c1908_wire_35_4, c1908_wire_35_5, c1908_wire_35_6});
fanout_n #(3, 0, 0) FANOUT_15 (c1908_wire_115, {c1908_wire_115_0, c1908_wire_115_1, c1908_wire_115_2});
fanout_n #(4, 0, 0) FANOUT_16 (c1908_wire_49, {c1908_wire_49_0, c1908_wire_49_1, c1908_wire_49_2, c1908_wire_49_3});
fanout_n #(4, 0, 0) FANOUT_17 (c1908_wire_121, {c1908_wire_121_0, c1908_wire_121_1, c1908_wire_121_2, c1908_wire_121_3});
fanout_n #(2, 0, 0) FANOUT_18 (c1908_wire_135, {c1908_wire_135_0, c1908_wire_135_1});
fanout_n #(5, 0, 0) FANOUT_19 (c1908_wire_125, {c1908_wire_125_0, c1908_wire_125_1, c1908_wire_125_2, c1908_wire_125_3, c1908_wire_125_4});
fanout_n #(3, 0, 0) FANOUT_20 (c1908_wire_140, {c1908_wire_140_0, c1908_wire_140_1, c1908_wire_140_2});
fanout_n #(6, 0, 0) FANOUT_21 (c1908_wire_30, {c1908_wire_30_0, c1908_wire_30_1, c1908_wire_30_2, c1908_wire_30_3, c1908_wire_30_4, c1908_wire_30_5});
fanout_n #(10, 0, 0) FANOUT_22 (c1908_wire_151, {c1908_wire_151_0, c1908_wire_151_1, c1908_wire_151_2, c1908_wire_151_3, c1908_wire_151_4, c1908_wire_151_5, c1908_wire_151_6, c1908_wire_151_7, c1908_wire_151_8, c1908_wire_151_9});
fanout_n #(10, 0, 0) FANOUT_23 (c1908_wire_155, {c1908_wire_155_0, c1908_wire_155_1, c1908_wire_155_2, c1908_wire_155_3, c1908_wire_155_4, c1908_wire_155_5, c1908_wire_155_6, c1908_wire_155_7, c1908_wire_155_8, c1908_wire_155_9});
fanout_n #(2, 0, 0) FANOUT_24 (c1908_wire_185, {c1908_wire_185_0, c1908_wire_185_1});
fanout_n #(10, 0, 0) FANOUT_25 (c1908_wire_156, {c1908_wire_156_0, c1908_wire_156_1, c1908_wire_156_2, c1908_wire_156_3, c1908_wire_156_4, c1908_wire_156_5, c1908_wire_156_6, c1908_wire_156_7, c1908_wire_156_8, c1908_wire_156_9});
fanout_n #(4, 0, 0) FANOUT_26 (c1908_wire_200, {c1908_wire_200_0, c1908_wire_200_1, c1908_wire_200_2, c1908_wire_200_3});
fanout_n #(5, 0, 0) FANOUT_27 (c1908_wire_211, {c1908_wire_211_0, c1908_wire_211_1, c1908_wire_211_2, c1908_wire_211_3, c1908_wire_211_4});
fanout_n #(7, 0, 0) FANOUT_28 (c1908_wire_67, {c1908_wire_67_0, c1908_wire_67_1, c1908_wire_67_2, c1908_wire_67_3, c1908_wire_67_4, c1908_wire_67_5, c1908_wire_67_6});
fanout_n #(10, 0, 0) FANOUT_29 (c1908_wire_157, {c1908_wire_157_0, c1908_wire_157_1, c1908_wire_157_2, c1908_wire_157_3, c1908_wire_157_4, c1908_wire_157_5, c1908_wire_157_6, c1908_wire_157_7, c1908_wire_157_8, c1908_wire_157_9});
fanout_n #(7, 0, 0) FANOUT_30 (c1908_wire_167, {c1908_wire_167_0, c1908_wire_167_1, c1908_wire_167_2, c1908_wire_167_3, c1908_wire_167_4, c1908_wire_167_5, c1908_wire_167_6});
fanout_n #(6, 0, 0) FANOUT_31 (c1908_wire_233, {c1908_wire_233_0, c1908_wire_233_1, c1908_wire_233_2, c1908_wire_233_3, c1908_wire_233_4, c1908_wire_233_5});
fanout_n #(2, 0, 0) FANOUT_32 (c1908_wire_56, {c1908_wire_56_0, c1908_wire_56_1});
fanout_n #(8, 0, 0) FANOUT_33 (c1908_wire_21, {c1908_wire_21_0, c1908_wire_21_1, c1908_wire_21_2, c1908_wire_21_3, c1908_wire_21_4, c1908_wire_21_5, c1908_wire_21_6, c1908_wire_21_7});
fanout_n #(5, 0, 0) FANOUT_34 (c1908_wire_241, {c1908_wire_241_0, c1908_wire_241_1, c1908_wire_241_2, c1908_wire_241_3, c1908_wire_241_4});
fanout_n #(6, 0, 0) FANOUT_35 (c1908_wire_22, {c1908_wire_22_0, c1908_wire_22_1, c1908_wire_22_2, c1908_wire_22_3, c1908_wire_22_4, c1908_wire_22_5});
fanout_n #(3, 0, 0) FANOUT_36 (c1908_wire_161, {c1908_wire_161_0, c1908_wire_161_1, c1908_wire_161_2});
fanout_n #(10, 0, 0) FANOUT_37 (c1908_wire_258, {c1908_wire_258_0, c1908_wire_258_1, c1908_wire_258_2, c1908_wire_258_3, c1908_wire_258_4, c1908_wire_258_5, c1908_wire_258_6, c1908_wire_258_7, c1908_wire_258_8, c1908_wire_258_9});
fanout_n #(7, 0, 0) FANOUT_38 (c1908_wire_70, {c1908_wire_70_0, c1908_wire_70_1, c1908_wire_70_2, c1908_wire_70_3, c1908_wire_70_4, c1908_wire_70_5, c1908_wire_70_6});
fanout_n #(7, 0, 0) FANOUT_39 (c1908_wire_218, {c1908_wire_218_0, c1908_wire_218_1, c1908_wire_218_2, c1908_wire_218_3, c1908_wire_218_4, c1908_wire_218_5, c1908_wire_218_6});
fanout_n #(10, 0, 0) FANOUT_40 (c1908_wire_277, {c1908_wire_277_0, c1908_wire_277_1, c1908_wire_277_2, c1908_wire_277_3, c1908_wire_277_4, c1908_wire_277_5, c1908_wire_277_6, c1908_wire_277_7, c1908_wire_277_8, c1908_wire_277_9});
fanout_n #(3, 0, 0) FANOUT_41 (c1908_wire_287, {c1908_wire_287_0, c1908_wire_287_1, c1908_wire_287_2});
fanout_n #(9, 0, 0) FANOUT_42 (c1908_wire_101, {c1908_wire_101_0, c1908_wire_101_1, c1908_wire_101_2, c1908_wire_101_3, c1908_wire_101_4, c1908_wire_101_5, c1908_wire_101_6, c1908_wire_101_7, c1908_wire_101_8});
fanout_n #(4, 0, 0) FANOUT_43 (c1908_wire_290, {c1908_wire_290_0, c1908_wire_290_1, c1908_wire_290_2, c1908_wire_290_3});
fanout_n #(6, 0, 0) FANOUT_44 (c1908_wire_291, {c1908_wire_291_0, c1908_wire_291_1, c1908_wire_291_2, c1908_wire_291_3, c1908_wire_291_4, c1908_wire_291_5});
fanout_n #(5, 0, 0) FANOUT_45 (c1908_wire_235, {c1908_wire_235_0, c1908_wire_235_1, c1908_wire_235_2, c1908_wire_235_3, c1908_wire_235_4});
fanout_n #(4, 0, 0) FANOUT_46 (c1908_wire_302, {c1908_wire_302_0, c1908_wire_302_1, c1908_wire_302_2, c1908_wire_302_3});
fanout_n #(2, 0, 0) FANOUT_47 (c1908_wire_137, {c1908_wire_137_0, c1908_wire_137_1});
fanout_n #(2, 0, 0) FANOUT_48 (c1908_wire_203, {c1908_wire_203_0, c1908_wire_203_1});
fanout_n #(4, 0, 0) FANOUT_49 (c1908_wire_318, {c1908_wire_318_0, c1908_wire_318_1, c1908_wire_318_2, c1908_wire_318_3});
fanout_n #(2, 0, 0) FANOUT_50 (c1908_wire_252, {c1908_wire_252_0, c1908_wire_252_1});
fanout_n #(5, 0, 0) FANOUT_51 (c1908_wire_197, {c1908_wire_197_0, c1908_wire_197_1, c1908_wire_197_2, c1908_wire_197_3, c1908_wire_197_4});
fanout_n #(2, 0, 0) FANOUT_52 (c1908_wire_79, {c1908_wire_79_0, c1908_wire_79_1});
fanout_n #(5, 0, 0) FANOUT_53 (c1908_wire_143, {c1908_wire_143_0, c1908_wire_143_1, c1908_wire_143_2, c1908_wire_143_3, c1908_wire_143_4});
fanout_n #(6, 0, 0) FANOUT_54 (c1908_wire_11, {c1908_wire_11_0, c1908_wire_11_1, c1908_wire_11_2, c1908_wire_11_3, c1908_wire_11_4, c1908_wire_11_5});
fanout_n #(2, 0, 0) FANOUT_55 (c1908_wire_408, {c1908_wire_408_0, c1908_wire_408_1});
fanout_n #(7, 0, 0) FANOUT_56 (c1908_wire_169, {c1908_wire_169_0, c1908_wire_169_1, c1908_wire_169_2, c1908_wire_169_3, c1908_wire_169_4, c1908_wire_169_5, c1908_wire_169_6});
fanout_n #(2, 0, 0) FANOUT_57 (c1908_wire_213, {c1908_wire_213_0, c1908_wire_213_1});
fanout_n #(3, 0, 0) FANOUT_58 (c1908_wire_85, {c1908_wire_85_0, c1908_wire_85_1, c1908_wire_85_2});
fanout_n #(6, 0, 0) FANOUT_59 (c1908_wire_52, {c1908_wire_52_0, c1908_wire_52_1, c1908_wire_52_2, c1908_wire_52_3, c1908_wire_52_4, c1908_wire_52_5});
fanout_n #(7, 0, 0) FANOUT_60 (c1908_wire_193, {c1908_wire_193_0, c1908_wire_193_1, c1908_wire_193_2, c1908_wire_193_3, c1908_wire_193_4, c1908_wire_193_5, c1908_wire_193_6});
fanout_n #(5, 0, 0) FANOUT_61 (c1908_wire_300, {c1908_wire_300_0, c1908_wire_300_1, c1908_wire_300_2, c1908_wire_300_3, c1908_wire_300_4});
fanout_n #(3, 0, 0) FANOUT_62 (c1908_wire_413, {c1908_wire_413_0, c1908_wire_413_1, c1908_wire_413_2});
fanout_n #(3, 0, 0) FANOUT_63 (c1908_wire_231, {c1908_wire_231_0, c1908_wire_231_1, c1908_wire_231_2});
fanout_n #(3, 0, 0) FANOUT_64 (c1908_wire_216, {c1908_wire_216_0, c1908_wire_216_1, c1908_wire_216_2});
fanout_n #(3, 0, 0) FANOUT_65 (c1908_wire_183, {c1908_wire_183_0, c1908_wire_183_1, c1908_wire_183_2});
fanout_n #(3, 0, 0) FANOUT_66 (c1908_wire_172, {c1908_wire_172_0, c1908_wire_172_1, c1908_wire_172_2});
fanout_n #(3, 0, 0) FANOUT_67 (c1908_wire_150, {c1908_wire_150_0, c1908_wire_150_1, c1908_wire_150_2});
fanout_n #(6, 0, 0) FANOUT_68 (c1908_wire_12, {c1908_wire_12_0, c1908_wire_12_1, c1908_wire_12_2, c1908_wire_12_3, c1908_wire_12_4, c1908_wire_12_5});
fanout_n #(3, 0, 0) FANOUT_69 (c1908_wire_387, {c1908_wire_387_0, c1908_wire_387_1, c1908_wire_387_2});
fanout_n #(21, 0, 0) FANOUT_70 (c1908_wire_96, {c1908_wire_96_0, c1908_wire_96_1, c1908_wire_96_2, c1908_wire_96_3, c1908_wire_96_4, c1908_wire_96_5, c1908_wire_96_6, c1908_wire_96_7, c1908_wire_96_8, c1908_wire_96_9, c1908_wire_96_10, c1908_wire_96_11, c1908_wire_96_12, c1908_wire_96_13, c1908_wire_96_14, c1908_wire_96_15, c1908_wire_96_16, c1908_wire_96_17, c1908_wire_96_18, c1908_wire_96_19, c1908_wire_96_20});
fanout_n #(3, 0, 0) FANOUT_71 (c1908_wire_361, {c1908_wire_361_0, c1908_wire_361_1, c1908_wire_361_2});
fanout_n #(6, 0, 0) FANOUT_72 (c1908_wire_365, {c1908_wire_365_0, c1908_wire_365_1, c1908_wire_365_2, c1908_wire_365_3, c1908_wire_365_4, c1908_wire_365_5});
fanout_n #(19, 0, 0) FANOUT_73 (c1908_wire_54, {c1908_wire_54_0, c1908_wire_54_1, c1908_wire_54_2, c1908_wire_54_3, c1908_wire_54_4, c1908_wire_54_5, c1908_wire_54_6, c1908_wire_54_7, c1908_wire_54_8, c1908_wire_54_9, c1908_wire_54_10, c1908_wire_54_11, c1908_wire_54_12, c1908_wire_54_13, c1908_wire_54_14, c1908_wire_54_15, c1908_wire_54_16, c1908_wire_54_17, c1908_wire_54_18});
fanout_n #(4, 0, 0) FANOUT_74 (c1908_wire_237, {c1908_wire_237_0, c1908_wire_237_1, c1908_wire_237_2, c1908_wire_237_3});
fanout_n #(7, 0, 0) FANOUT_75 (c1908_wire_239, {c1908_wire_239_0, c1908_wire_239_1, c1908_wire_239_2, c1908_wire_239_3, c1908_wire_239_4, c1908_wire_239_5, c1908_wire_239_6});
fanout_n #(4, 0, 0) FANOUT_76 (c1908_wire_303, {c1908_wire_303_0, c1908_wire_303_1, c1908_wire_303_2, c1908_wire_303_3});
fanout_n #(6, 0, 0) FANOUT_77 (c1908_wire_43, {c1908_wire_43_0, c1908_wire_43_1, c1908_wire_43_2, c1908_wire_43_3, c1908_wire_43_4, c1908_wire_43_5});
fanout_n #(5, 0, 0) FANOUT_78 (c1908_wire_163, {c1908_wire_163_0, c1908_wire_163_1, c1908_wire_163_2, c1908_wire_163_3, c1908_wire_163_4});
fanout_n #(6, 0, 0) FANOUT_79 (c1908_wire_41, {c1908_wire_41_0, c1908_wire_41_1, c1908_wire_41_2, c1908_wire_41_3, c1908_wire_41_4, c1908_wire_41_5});
fanout_n #(6, 0, 0) FANOUT_80 (c1908_wire_42, {c1908_wire_42_0, c1908_wire_42_1, c1908_wire_42_2, c1908_wire_42_3, c1908_wire_42_4, c1908_wire_42_5});
fanout_n #(2, 0, 0) FANOUT_81 (c1908_wire_36, {c1908_wire_36_0, c1908_wire_36_1});
fanout_n #(5, 0, 0) FANOUT_82 (c1908_wire_106, {c1908_wire_106_0, c1908_wire_106_1, c1908_wire_106_2, c1908_wire_106_3, c1908_wire_106_4});
fanout_n #(2, 0, 0) FANOUT_83 (c1908_wire_111, {c1908_wire_111_0, c1908_wire_111_1});
fanout_n #(3, 0, 0) FANOUT_84 (c1908_wire_265, {c1908_wire_265_0, c1908_wire_265_1, c1908_wire_265_2});
fanout_n #(3, 0, 0) FANOUT_85 (c1908_wire_268, {c1908_wire_268_0, c1908_wire_268_1, c1908_wire_268_2});
fanout_n #(8, 0, 0) FANOUT_86 (c1908_wire_279, {c1908_wire_279_0, c1908_wire_279_1, c1908_wire_279_2, c1908_wire_279_3, c1908_wire_279_4, c1908_wire_279_5, c1908_wire_279_6, c1908_wire_279_7});
fanout_n #(7, 0, 0) FANOUT_87 (c1908_wire_15, {c1908_wire_15_0, c1908_wire_15_1, c1908_wire_15_2, c1908_wire_15_3, c1908_wire_15_4, c1908_wire_15_5, c1908_wire_15_6});
fanout_n #(2, 0, 0) FANOUT_88 (c1908_wire_112, {c1908_wire_112_0, c1908_wire_112_1});
fanout_n #(4, 0, 0) FANOUT_89 (c1908_wire_87, {c1908_wire_87_0, c1908_wire_87_1, c1908_wire_87_2, c1908_wire_87_3});
fanout_n #(4, 0, 0) FANOUT_90 (c1908_wire_88, {c1908_wire_88_0, c1908_wire_88_1, c1908_wire_88_2, c1908_wire_88_3});
fanout_n #(2, 0, 0) FANOUT_91 (c1908_wire_76, {c1908_wire_76_0, c1908_wire_76_1});
fanout_n #(2, 0, 0) FANOUT_92 (c1908_wire_77, {c1908_wire_77_0, c1908_wire_77_1});


bufg #(0, 0) BUF_1 (c1908_wire_1, G1_net_0);
bufg #(0, 0) BUF_2 (c1908_wire_2, G10_net_0);
and_n #(2, 0, 0) AND_1 (c1908_wire_3, {c1908_wire_4_0, c1908_wire_5_0});
and_n #(2, 0, 0) AND_2 (c1908_wire_6, {c1908_wire_4_1, c1908_wire_7});
or_n #(2, 0, 0) OR_1 (c1908_wire_4, {c1908_wire_8, c1908_wire_9});
xor_n #(2, 0, 0) XOR_1 (c1908_wire_10, {c1908_wire_11_0, c1908_wire_12_0});
and_n #(2, 0, 0) AND_3 (c1908_wire_8, {c1908_wire_10, c1908_wire_1_0});
nor_n #(2, 0, 0) NOR_1 (c1908_wire_9, {c1908_wire_1_1, c1908_wire_13});
xor_n #(2, 0, 0) XOR_2 (c1908_wire_13, {c1908_wire_11_1, c1908_wire_12_1});
xor_n #(2, 0, 0) XOR_3 (c1908_wire_14, {c1908_wire_5_1, c1908_wire_15_0});
and_n #(2, 0, 0) AND_4 (c1908_wire_16, {c1908_wire_5_2, c1908_wire_17_0});
or_n #(2, 0, 0) OR_2 (c1908_wire_5, {c1908_wire_18, c1908_wire_19});
xor_n #(2, 0, 0) XOR_4 (c1908_wire_20, {c1908_wire_21_0, c1908_wire_22_0});
and_n #(2, 0, 0) AND_5 (c1908_wire_18, {c1908_wire_20, c1908_wire_2_0});
nor_n #(2, 0, 0) NOR_2 (c1908_wire_19, {c1908_wire_2_1, c1908_wire_23});
xor_n #(2, 0, 0) XOR_5 (c1908_wire_23, {c1908_wire_21_1, c1908_wire_22_1});
and_n #(2, 0, 0) AND_6 (c1908_wire_24, {c1908_wire_17_1, c1908_wire_25});
or_n #(2, 0, 0) OR_3 (c1908_wire_17, {c1908_wire_26, c1908_wire_27});
xor_n #(2, 0, 0) XOR_6 (c1908_wire_28, {c1908_wire_29_0, c1908_wire_30_0});
and_n #(2, 0, 0) AND_7 (c1908_wire_26, {c1908_wire_28, c1908_wire_31_0});
nor_n #(2, 0, 0) NOR_3 (c1908_wire_27, {c1908_wire_31_1, c1908_wire_32});
xor_n #(2, 0, 0) XOR_7 (c1908_wire_32, {c1908_wire_29_1, c1908_wire_30_1});
and_n #(2, 0, 0) AND_8 (c1908_wire_33, {c1908_wire_34_0, c1908_wire_35_0});
xor_n #(2, 0, 0) XOR_8 (c1908_wire_7, {c1908_wire_34_1, c1908_wire_36_0});
xor_n #(2, 0, 0) XOR_9 (c1908_wire_37, {c1908_wire_34_2, c1908_wire_36_1});
or_n #(2, 0, 0) OR_4 (c1908_wire_34, {c1908_wire_38, c1908_wire_39});
xor_n #(2, 0, 0) XOR_10 (c1908_wire_40, {c1908_wire_41_0, c1908_wire_42_0});
and_n #(2, 0, 0) AND_9 (c1908_wire_38, {c1908_wire_40, c1908_wire_43_0});
nor_n #(2, 0, 0) NOR_4 (c1908_wire_39, {c1908_wire_43_1, c1908_wire_44});
xor_n #(2, 0, 0) XOR_11 (c1908_wire_44, {c1908_wire_41_1, c1908_wire_42_1});
or_n #(2, 0, 0) OR_5 (c1908_wire_45, {c1908_wire_46, c1908_wire_47});
and_n #(2, 0, 0) AND_10 (c1908_wire_48, {c1908_wire_45_0, c1908_wire_49_0});
and_n #(2, 0, 0) AND_11 (c1908_wire_50, {c1908_wire_45_1, c1908_wire_49_1});
notg #(0, 0) NOT_1 (c1908_wire_51, c1908_wire_52_0);
or_n #(2, 0, 0) OR_6 (c1908_wire_53, {c1908_wire_51, c1908_wire_54_0});
notg #(0, 0) NOT_2 (c1908_wire_55, c1908_wire_56_0);
and_n #(2, 0, 0) AND_12 (c1908_wire_47, {c1908_wire_55, c1908_wire_53});
and_n #(2, 0, 0) AND_13 (c1908_wire_57, {c1908_wire_52_1, c1908_wire_56_1});
and_n #(2, 0, 0) AND_14 (c1908_wire_46, {c1908_wire_57, c1908_wire_58});
notg #(0, 0) NOT_3 (c1908_wire_58, c1908_wire_54_1);
and_n #(2, 0, 0) AND_15 (c1908_wire_59, {c1908_wire_60_0, c1908_wire_61});
and_n #(2, 0, 0) AND_16 (c1908_wire_62, {c1908_wire_60_1, c1908_wire_63});
or_n #(2, 0, 0) OR_7 (c1908_wire_60, {c1908_wire_64, c1908_wire_65});
xor_n #(2, 0, 0) XOR_12 (c1908_wire_66, {c1908_wire_22_2, c1908_wire_15_1});
and_n #(2, 0, 0) AND_17 (c1908_wire_64, {c1908_wire_66, c1908_wire_67_0});
nor_n #(2, 0, 0) NOR_5 (c1908_wire_65, {c1908_wire_67_1, c1908_wire_68});
xor_n #(2, 0, 0) XOR_13 (c1908_wire_68, {c1908_wire_22_3, c1908_wire_15_2});
and_n #(2, 0, 0) AND_18 (c1908_wire_69, {c1908_wire_2_2, c1908_wire_70_0});
and_n #(2, 0, 0) AND_19 (c1908_wire_71, {c1908_wire_2_3, c1908_wire_72});
and_n #(2, 0, 0) AND_20 (c1908_wire_73, {c1908_wire_2_4, c1908_wire_74});
bufg #(0, 0) BUF_3 (c1908_wire_31, G11_net_0);
xor_n #(2, 0, 0) XOR_14 (c1908_wire_75, {c1908_wire_76_0, c1908_wire_77_0});
and_n #(2, 0, 0) AND_21 (c1908_wire_78, {c1908_wire_75, c1908_wire_79_0});
nor_n #(2, 0, 0) NOR_6 (c1908_wire_80, {c1908_wire_79_1, c1908_wire_81});
xor_n #(2, 0, 0) XOR_15 (c1908_wire_81, {c1908_wire_76_1, c1908_wire_77_1});
or_n #(2, 0, 0) OR_8 (c1908_wire_82, {c1908_wire_78, c1908_wire_80});
notg #(0, 0) NOT_4 (c1908_wire_83, c1908_wire_14_0);
and_n #(2, 0, 0) AND_22 (c1908_wire_84, {c1908_wire_14_1, c1908_wire_85_0});
and_n #(2, 0, 0) AND_23 (c1908_wire_86, {c1908_wire_87_0, c1908_wire_88_0});
or_n #(2, 0, 0) OR_9 (c1908_wire_61, {c1908_wire_86, c1908_wire_89});
nor_n #(2, 0, 0) NOR_7 (c1908_wire_89, {c1908_wire_87_1, c1908_wire_88_1});
or_n #(2, 0, 0) OR_10 (c1908_wire_90, {c1908_wire_91, c1908_wire_92});
or_n #(2, 0, 0) OR_11 (c1908_wire_93, {c1908_wire_59, c1908_wire_94});
nor_n #(2, 0, 0) NOR_8 (c1908_wire_94, {c1908_wire_90, c1908_wire_60_2});
and_n #(2, 0, 0) AND_24 (c1908_wire_91, {c1908_wire_87_2, c1908_wire_88_2});
nor_n #(2, 0, 0) NOR_9 (c1908_wire_92, {c1908_wire_87_3, c1908_wire_88_3});
or_n #(2, 0, 0) OR_12 (c1908_wire_95, {c1908_wire_82_0, c1908_wire_96_0});
notg #(0, 0) NOT_5 (c1908_wire_97, c1908_wire_82_1);
xor_n #(2, 0, 0) XOR_16 (c1908_wire_98, {c1908_wire_82_2, c1908_wire_99});
and_n #(2, 0, 0) AND_25 (c1908_wire_100, {c1908_wire_31_2, c1908_wire_101_0});
and_n #(2, 0, 0) AND_26 (c1908_wire_102, {c1908_wire_31_3, c1908_wire_103});
bufg #(0, 0) BUF_4 (c1908_wire_29, G12_net_0);
or_n #(2, 0, 0) OR_13 (c1908_wire_35, {c1908_wire_16, c1908_wire_104});
xor_n #(2, 0, 0) XOR_17 (c1908_wire_105, {c1908_wire_35_1, c1908_wire_106_0});
xor_n #(2, 0, 0) XOR_18 (c1908_wire_107, {c1908_wire_35_2, c1908_wire_106_1});
xor_n #(2, 0, 0) XOR_19 (c1908_wire_108, {c1908_wire_35_3, c1908_wire_106_2});
xor_n #(2, 0, 0) XOR_20 (c1908_wire_109, {c1908_wire_35_4, c1908_wire_106_3});
xor_n #(2, 0, 0) XOR_21 (c1908_wire_110, {c1908_wire_35_5, c1908_wire_106_4});
nor_n #(2, 0, 0) NOR_10 (c1908_wire_104, {c1908_wire_5_3, c1908_wire_17_2});
xor_n #(2, 0, 0) XOR_22 (c1908_wire_63, {c1908_wire_111_0, c1908_wire_112_0});
nor_n #(2, 0, 0) NOR_11 (c1908_wire_113, {c1908_wire_60_3, c1908_wire_114});
xor_n #(2, 0, 0) XOR_23 (c1908_wire_114, {c1908_wire_111_1, c1908_wire_112_1});
or_n #(2, 0, 0) OR_14 (c1908_wire_115, {c1908_wire_62, c1908_wire_113});
or_n #(2, 0, 0) OR_15 (c1908_wire_116, {c1908_wire_93_0, c1908_wire_96_1});
notg #(0, 0) NOT_6 (c1908_wire_117, c1908_wire_93_1);
xor_n #(2, 0, 0) XOR_24 (c1908_wire_118, {c1908_wire_93_2, c1908_wire_119});
or_n #(2, 0, 0) OR_16 (c1908_wire_49, {c1908_wire_3, c1908_wire_120});
nor_n #(2, 0, 0) NOR_12 (c1908_wire_120, {c1908_wire_4_2, c1908_wire_5_4});
or_n #(2, 0, 0) OR_17 (c1908_wire_121, {c1908_wire_122, c1908_wire_123});
and_n #(2, 0, 0) AND_27 (c1908_wire_124, {c1908_wire_121_0, c1908_wire_125_0});
and_n #(2, 0, 0) AND_28 (c1908_wire_126, {c1908_wire_121_1, c1908_wire_127});
notg #(0, 0) NOT_7 (c1908_wire_128, c1908_wire_85_1);
or_n #(2, 0, 0) OR_18 (c1908_wire_129, {c1908_wire_128, c1908_wire_54_2});
and_n #(2, 0, 0) AND_29 (c1908_wire_123, {c1908_wire_83, c1908_wire_129});
and_n #(2, 0, 0) AND_30 (c1908_wire_122, {c1908_wire_84, c1908_wire_130});
notg #(0, 0) NOT_8 (c1908_wire_130, c1908_wire_54_3);
xor_n #(2, 0, 0) XOR_25 (c1908_wire_131, {c1908_wire_115_0, c1908_wire_132});
and_n #(2, 0, 0) AND_31 (c1908_wire_133, {c1908_wire_115_1, c1908_wire_134});
and_n #(2, 0, 0) AND_32 (c1908_wire_135, {c1908_wire_125_1, c1908_wire_136});
xor_n #(2, 0, 0) XOR_26 (c1908_wire_127, {c1908_wire_125_2, c1908_wire_137_0});
xor_n #(2, 0, 0) XOR_27 (c1908_wire_138, {c1908_wire_125_3, c1908_wire_137_1});
or_n #(2, 0, 0) OR_19 (c1908_wire_125, {c1908_wire_6, c1908_wire_139});
nor_n #(2, 0, 0) NOR_13 (c1908_wire_139, {c1908_wire_4_3, c1908_wire_37});
or_n #(2, 0, 0) OR_20 (c1908_wire_140, {c1908_wire_33, c1908_wire_141});
xor_n #(2, 0, 0) XOR_28 (c1908_wire_142, {c1908_wire_140_0, c1908_wire_143_0});
and_n #(2, 0, 0) AND_33 (c1908_wire_144, {c1908_wire_140_1, c1908_wire_145});
nor_n #(2, 0, 0) NOR_14 (c1908_wire_141, {c1908_wire_35_6, c1908_wire_34_3});
and_n #(2, 0, 0) AND_34 (c1908_wire_146, {c1908_wire_29_2, c1908_wire_101_1});
xor_n #(2, 0, 0) XOR_29 (c1908_wire_74, {c1908_wire_29_3, c1908_wire_21_2});
xor_n #(2, 0, 0) XOR_30 (c1908_wire_147, {c1908_wire_29_4, c1908_wire_21_3});
bufg #(0, 0) BUF_5 (c1908_wire_30, G13_net_0);
and_n #(2, 0, 0) AND_35 (c1908_wire_148, {c1908_wire_135_0, c1908_wire_149});
or_n #(2, 0, 0) OR_21 (c1908_wire_136, {c1908_wire_150_0, c1908_wire_54_4});
or_n #(2, 0, 0) OR_22 (c1908_wire_151, {c1908_wire_152, c1908_wire_153});
and_n #(4, 0, 0) AND_36 (c1908_wire_154, {c1908_wire_151_0, c1908_wire_155_0, c1908_wire_156_0, c1908_wire_157_0});
and_n #(4, 0, 0) AND_37 (c1908_wire_158, {c1908_wire_151_1, c1908_wire_155_1, c1908_wire_156_1, c1908_wire_157_1});
and_n #(4, 0, 0) AND_38 (c1908_wire_159, {c1908_wire_151_2, c1908_wire_155_2, c1908_wire_156_2, c1908_wire_157_2});
and_n #(4, 0, 0) AND_39 (c1908_wire_160, {c1908_wire_151_3, c1908_wire_156_3, c1908_wire_157_3, c1908_wire_161_0});
and_n #(4, 0, 0) AND_40 (c1908_wire_162, {c1908_wire_151_4, c1908_wire_156_4, c1908_wire_161_1, c1908_wire_163_0});
and_n #(2, 0, 0) AND_41 (c1908_wire_164, {c1908_wire_151_5, c1908_wire_155_3});
and_n #(2, 0, 0) AND_42 (c1908_wire_165, {c1908_wire_151_6, c1908_wire_155_4});
and_n #(2, 0, 0) AND_43 (c1908_wire_166, {c1908_wire_151_7, c1908_wire_167_0});
and_n #(8, 0, 0) AND_44 (c1908_wire_168, {c1908_wire_151_8, c1908_wire_155_5, c1908_wire_156_5, c1908_wire_157_4, c1908_wire_167_1, c1908_wire_161_2, c1908_wire_163_1, c1908_wire_169_0});
and_n #(4, 0, 0) AND_45 (c1908_wire_170, {c1908_wire_151_9, c1908_wire_155_6, c1908_wire_156_6, c1908_wire_157_5});
and_n #(2, 0, 0) AND_46 (c1908_wire_152, {c1908_wire_95, c1908_wire_171});
notg #(0, 0) NOT_9 (c1908_wire_171, c1908_wire_172_0);
and_n #(3, 0, 0) AND_47 (c1908_wire_153, {c1908_wire_97, c1908_wire_173, c1908_wire_172_1});
notg #(0, 0) NOT_10 (c1908_wire_173, c1908_wire_96_2);
or_n #(2, 0, 0) OR_23 (c1908_wire_155, {c1908_wire_174, c1908_wire_175});
and_n #(3, 0, 0) AND_48 (c1908_wire_176, {c1908_wire_155_7, c1908_wire_177, c1908_wire_178});
and_n #(2, 0, 0) AND_49 (c1908_wire_179, {c1908_wire_155_8, c1908_wire_157_6});
and_n #(2, 0, 0) AND_50 (c1908_wire_180, {c1908_wire_155_9, c1908_wire_181});
and_n #(2, 0, 0) AND_51 (c1908_wire_174, {c1908_wire_116, c1908_wire_182});
notg #(0, 0) NOT_11 (c1908_wire_182, c1908_wire_183_0);
and_n #(3, 0, 0) AND_52 (c1908_wire_175, {c1908_wire_117, c1908_wire_184, c1908_wire_183_1});
notg #(0, 0) NOT_12 (c1908_wire_184, c1908_wire_96_3);
and_n #(2, 0, 0) AND_53 (c1908_wire_185, {c1908_wire_142, c1908_wire_186});
notg #(0, 0) NOT_13 (c1908_wire_186, c1908_wire_96_4);
and_n #(4, 0, 0) AND_54 (c1908_wire_187, {c1908_wire_156_7, c1908_wire_157_7, c1908_wire_167_2, c1908_wire_169_1});
and_n #(4, 0, 0) AND_55 (c1908_wire_188, {c1908_wire_156_8, c1908_wire_157_8, c1908_wire_167_3, c1908_wire_169_2});
and_n #(4, 0, 0) AND_56 (c1908_wire_189, {c1908_wire_156_9, c1908_wire_157_9, c1908_wire_163_2, c1908_wire_169_3});
or_n #(3, 0, 0) OR_24 (c1908_wire_156, {c1908_wire_190, c1908_wire_133, c1908_wire_191});
nor_n #(2, 0, 0) NOR_15 (c1908_wire_192, {c1908_wire_193_0, c1908_wire_96_5});
nor_n #(2, 0, 0) NOR_16 (c1908_wire_194, {c1908_wire_115_2, c1908_wire_96_6});
and_n #(2, 0, 0) AND_57 (c1908_wire_190, {c1908_wire_194, c1908_wire_195});
or_n #(2, 0, 0) OR_25 (c1908_wire_134, {c1908_wire_196, c1908_wire_192});
notg #(0, 0) NOT_14 (c1908_wire_196, c1908_wire_197_0);
notg #(0, 0) NOT_15 (c1908_wire_198, c1908_wire_197_1);
and_n #(2, 0, 0) AND_58 (c1908_wire_191, {c1908_wire_198, c1908_wire_96_7});
and_n #(2, 0, 0) AND_59 (c1908_wire_195, {c1908_wire_197_2, c1908_wire_193_1});
or_n #(2, 0, 0) OR_26 (c1908_wire_199, {c1908_wire_200_0, c1908_wire_96_8});
notg #(0, 0) NOT_16 (c1908_wire_201, c1908_wire_200_1);
and_n #(2, 0, 0) AND_60 (c1908_wire_202, {c1908_wire_200_2, c1908_wire_203_0});
or_n #(2, 0, 0) OR_27 (c1908_wire_200, {c1908_wire_24, c1908_wire_204});
or_n #(2, 0, 0) OR_28 (c1908_wire_25, {c1908_wire_48, c1908_wire_205});
or_n #(2, 0, 0) OR_29 (c1908_wire_206, {c1908_wire_50, c1908_wire_207});
nor_n #(2, 0, 0) NOR_17 (c1908_wire_204, {c1908_wire_206, c1908_wire_17_3});
nor_n #(2, 0, 0) NOR_18 (c1908_wire_205, {c1908_wire_45_2, c1908_wire_49_2});
nor_n #(2, 0, 0) NOR_19 (c1908_wire_207, {c1908_wire_45_3, c1908_wire_49_3});
or_n #(2, 0, 0) OR_30 (c1908_wire_208, {c1908_wire_124, c1908_wire_209});
nor_n #(2, 0, 0) NOR_20 (c1908_wire_209, {c1908_wire_121_2, c1908_wire_125_4});
notg #(0, 0) NOT_17 (c1908_wire_210, c1908_wire_96_9);
and_n #(2, 0, 0) AND_61 (c1908_wire_211, {c1908_wire_210, c1908_wire_208});
and_n #(2, 0, 0) AND_62 (c1908_wire_212, {c1908_wire_30_2, c1908_wire_213_0});
and_n #(2, 0, 0) AND_63 (c1908_wire_214, {c1908_wire_30_3, c1908_wire_101_2});
bufg #(0, 0) BUF_6 (c1908_wire_67, G14_net_0);
and_n #(2, 0, 0) AND_64 (c1908_wire_215, {c1908_wire_185_0, c1908_wire_216_0});
xor_n #(2, 0, 0) XOR_31 (c1908_wire_217, {c1908_wire_211_0, c1908_wire_218_0});
and_n #(2, 0, 0) AND_65 (c1908_wire_219, {c1908_wire_211_1, c1908_wire_218_1});
notg #(0, 0) NOT_18 (c1908_wire_220, c1908_wire_211_2);
and_n #(2, 0, 0) AND_66 (c1908_wire_221, {c1908_wire_211_3, c1908_wire_218_2});
or_n #(2, 0, 0) OR_31 (c1908_wire_157, {c1908_wire_215, c1908_wire_222});
nor_n #(2, 0, 0) NOR_21 (c1908_wire_222, {c1908_wire_185_1, c1908_wire_216_1});
notg #(0, 0) NOT_19 (c1908_wire_223, c1908_wire_167_4);
or_n #(2, 0, 0) OR_32 (c1908_wire_167, {c1908_wire_224, c1908_wire_225});
and_n #(3, 0, 0) AND_67 (c1908_wire_226, {c1908_wire_167_5, c1908_wire_227, c1908_wire_228});
and_n #(2, 0, 0) AND_68 (c1908_wire_229, {c1908_wire_167_6, c1908_wire_169_4});
and_n #(2, 0, 0) AND_69 (c1908_wire_224, {c1908_wire_199, c1908_wire_230});
notg #(0, 0) NOT_20 (c1908_wire_230, c1908_wire_231_0);
and_n #(3, 0, 0) AND_70 (c1908_wire_225, {c1908_wire_201, c1908_wire_232, c1908_wire_231_1});
notg #(0, 0) NOT_21 (c1908_wire_232, c1908_wire_96_10);
and_n #(3, 0, 0) AND_71 (c1908_wire_233, {c1908_wire_217, c1908_wire_234, c1908_wire_235_0});
notg #(0, 0) NOT_22 (c1908_wire_181, c1908_wire_233_0);
notg #(0, 0) NOT_23 (c1908_wire_236, c1908_wire_233_1);
notg #(0, 0) NOT_24 (c1908_wire_234, c1908_wire_237_0);
and_n #(2, 0, 0) AND_72 (c1908_wire_238, {c1908_wire_67_2, c1908_wire_15_3});
xor_n #(2, 0, 0) XOR_32 (c1908_wire_56, {c1908_wire_67_3, c1908_wire_239_0});
and_n #(2, 0, 0) AND_73 (c1908_wire_240, {c1908_wire_67_4, c1908_wire_101_3});
bufg #(0, 0) BUF_7 (c1908_wire_21, G15_net_0);
and_n #(2, 0, 0) AND_74 (c1908_wire_241, {c1908_wire_223, c1908_wire_169_5});
notg #(0, 0) NOT_25 (c1908_wire_177, c1908_wire_241_0);
notg #(0, 0) NOT_26 (c1908_wire_242, c1908_wire_241_1);
notg #(0, 0) NOT_27 (c1908_wire_243, c1908_wire_241_2);
and_n #(2, 0, 0) AND_75 (c1908_wire_244, {c1908_wire_154, c1908_wire_226});
notg #(0, 0) NOT_28 (c1908_wire_245, c1908_wire_244);
nor_n #(2, 0, 0) NOR_22 (c1908_wire_246, {c1908_wire_235_1, c1908_wire_237_1});
and_n #(2, 0, 0) AND_76 (c1908_wire_247, {c1908_wire_246, c1908_wire_221});
or_n #(2, 0, 0) OR_33 (c1908_wire_248, {c1908_wire_249, c1908_wire_237_2});
and_n #(2, 0, 0) AND_77 (c1908_wire_250, {c1908_wire_248, c1908_wire_220});
or_n #(2, 0, 0) OR_34 (c1908_wire_227, {c1908_wire_247, c1908_wire_250});
nor_n #(2, 0, 0) NOR_23 (c1908_wire_249, {c1908_wire_218_3, c1908_wire_235_2});
notg #(0, 0) NOT_29 (c1908_wire_228, c1908_wire_169_6);
and_n #(2, 0, 0) AND_78 (c1908_wire_251, {c1908_wire_21_4, c1908_wire_70_1});
xor_n #(2, 0, 0) XOR_33 (c1908_wire_103, {c1908_wire_21_5, c1908_wire_252_0});
xor_n #(2, 0, 0) XOR_34 (c1908_wire_253, {c1908_wire_21_6, c1908_wire_252_1});
bufg #(0, 0) BUF_8 (c1908_wire_22, G16_net_0);
and_n #(3, 0, 0) AND_79 (c1908_wire_161, {c1908_wire_254, c1908_wire_255, c1908_wire_235_3});
or_n #(2, 0, 0) OR_35 (c1908_wire_255, {c1908_wire_219, c1908_wire_256});
nor_n #(2, 0, 0) NOR_24 (c1908_wire_256, {c1908_wire_211_4, c1908_wire_218_4});
notg #(0, 0) NOT_30 (c1908_wire_254, c1908_wire_237_3);
and_n #(2, 0, 0) AND_80 (c1908_wire_257, {c1908_wire_258_0, c1908_wire_1_2});
and_n #(2, 0, 0) AND_81 (c1908_wire_259, {c1908_wire_258_1, c1908_wire_11_2});
and_n #(2, 0, 0) AND_82 (c1908_wire_260, {c1908_wire_258_2, c1908_wire_12_2});
and_n #(2, 0, 0) AND_83 (c1908_wire_261, {c1908_wire_258_3, c1908_wire_239_1});
and_n #(2, 0, 0) AND_84 (c1908_wire_258, {c1908_wire_158, c1908_wire_262});
notg #(0, 0) NOT_31 (c1908_wire_263, c1908_wire_258_4);
notg #(0, 0) NOT_32 (c1908_wire_264, c1908_wire_258_5);
nor_n #(3, 0, 0) NOR_25 (c1908_wire_262, {c1908_wire_233_2, c1908_wire_241_3, c1908_wire_265_0});
and_n #(2, 0, 0) AND_85 (c1908_wire_266, {c1908_wire_70_2, c1908_wire_22_4});
and_n #(2, 0, 0) AND_86 (c1908_wire_70, {c1908_wire_159, c1908_wire_267});
nor_n #(3, 0, 0) NOR_26 (c1908_wire_267, {c1908_wire_233_3, c1908_wire_241_4, c1908_wire_268_0});
bufg #(0, 0) BUF_9 (c1908_wire_218, G17_net_0);
and_n #(2, 0, 0) AND_87 (c1908_wire_269, {c1908_wire_189, c1908_wire_270});
notg #(0, 0) NOT_33 (c1908_wire_271, c1908_wire_269);
and_n #(2, 0, 0) AND_88 (c1908_wire_270, {c1908_wire_166, c1908_wire_180});
and_n #(2, 0, 0) AND_89 (c1908_wire_272, {c1908_wire_162, c1908_wire_273});
notg #(0, 0) NOT_34 (c1908_wire_274, c1908_wire_272);
and_n #(2, 0, 0) AND_90 (c1908_wire_273, {c1908_wire_179, c1908_wire_242});
notg #(0, 0) NOT_35 (c1908_wire_275, c1908_wire_168);
and_n #(2, 0, 0) AND_91 (c1908_wire_276, {c1908_wire_277_0, c1908_wire_43_2});
and_n #(2, 0, 0) AND_92 (c1908_wire_278, {c1908_wire_277_1, c1908_wire_279_0});
and_n #(2, 0, 0) AND_93 (c1908_wire_280, {c1908_wire_277_2, c1908_wire_41_2});
and_n #(2, 0, 0) AND_94 (c1908_wire_281, {c1908_wire_277_3, c1908_wire_42_2});
and_n #(2, 0, 0) AND_95 (c1908_wire_277, {c1908_wire_187, c1908_wire_282});
notg #(0, 0) NOT_36 (c1908_wire_283, c1908_wire_277_4);
notg #(0, 0) NOT_37 (c1908_wire_284, c1908_wire_277_5);
and_n #(2, 0, 0) AND_96 (c1908_wire_282, {c1908_wire_164, c1908_wire_285});
nor_n #(2, 0, 0) NOR_27 (c1908_wire_285, {c1908_wire_233_4, c1908_wire_265_1});
and_n #(2, 0, 0) AND_97 (c1908_wire_286, {c1908_wire_287_0, c1908_wire_15_4});
and_n #(2, 0, 0) AND_98 (c1908_wire_287, {c1908_wire_188, c1908_wire_288});
and_n #(2, 0, 0) AND_99 (c1908_wire_288, {c1908_wire_165, c1908_wire_289});
nor_n #(2, 0, 0) NOR_28 (c1908_wire_289, {c1908_wire_233_5, c1908_wire_268_1});
and_n #(2, 0, 0) AND_100 (c1908_wire_101, {c1908_wire_160, c1908_wire_176});
notg #(0, 0) NOT_38 (c1908_wire_178, c1908_wire_268_2);
nor_n #(3, 0, 0) NOR_29 (c1908_wire_290, {c1908_wire_70_3, c1908_wire_287_1, c1908_wire_101_4});
and_n #(3, 0, 0) AND_101 (c1908_wire_291, {c1908_wire_290_0, c1908_wire_263, c1908_wire_283});
and_n #(6, 0, 0) AND_102 (c1908_wire_292, {c1908_wire_290_1, c1908_wire_271, c1908_wire_264, c1908_wire_274, c1908_wire_284, c1908_wire_275});
notg #(0, 0) NOT_39 (c1908_wire_293, c1908_wire_290_2);
and_n #(2, 0, 0) AND_103 (c1908_wire_294, {c1908_wire_290_3, c1908_wire_295});
and_n #(3, 0, 0) AND_104 (c1908_wire_296, {c1908_wire_218_5, c1908_wire_297, c1908_wire_298});
and_n #(2, 0, 0) AND_105 (c1908_wire_299, {c1908_wire_218_6, c1908_wire_300_0});
bufg #(0, 0) BUF_10 (c1908_wire_235, G18_net_0);
and_n #(2, 0, 0) AND_106 (c1908_wire_301, {c1908_wire_302_0, c1908_wire_303_0});
and_n #(2, 0, 0) AND_107 (c1908_wire_304, {c1908_wire_302_1, c1908_wire_303_1});
and_n #(2, 0, 0) AND_108 (c1908_wire_302, {c1908_wire_170, c1908_wire_305});
or_n #(2, 0, 0) OR_36 (c1908_wire_306, {c1908_wire_229, c1908_wire_243});
and_n #(3, 0, 0) AND_109 (c1908_wire_305, {c1908_wire_236, c1908_wire_306, c1908_wire_307});
nor_n #(2, 0, 0) NOR_30 (c1908_wire_307, {c1908_wire_54_5, c1908_wire_265_2});
notg #(0, 0) NOT_40 (c1908_wire_308, c1908_wire_291_0);
notg #(0, 0) NOT_41 (c1908_wire_309, c1908_wire_291_1);
notg #(0, 0) NOT_42 (c1908_wire_310, c1908_wire_291_2);
notg #(0, 0) NOT_43 (c1908_wire_311, c1908_wire_291_3);
and_n #(2, 0, 0) AND_110 (c1908_wire_137, {c1908_wire_299, c1908_wire_312});
nor_n #(2, 0, 0) NOR_31 (c1908_wire_312, {c1908_wire_96_11, c1908_wire_291_4});
and_n #(3, 0, 0) AND_111 (c1908_wire_203, {c1908_wire_313, c1908_wire_308, c1908_wire_231_2});
notg #(0, 0) NOT_44 (c1908_wire_313, c1908_wire_96_12);
and_n #(3, 0, 0) AND_112 (c1908_wire_119, {c1908_wire_314, c1908_wire_309, c1908_wire_183_2});
notg #(0, 0) NOT_45 (c1908_wire_314, c1908_wire_96_13);
and_n #(3, 0, 0) AND_113 (c1908_wire_99, {c1908_wire_315, c1908_wire_310, c1908_wire_172_2});
notg #(0, 0) NOT_46 (c1908_wire_315, c1908_wire_96_14);
and_n #(2, 0, 0) AND_114 (c1908_wire_132, {c1908_wire_316, c1908_wire_317});
and_n #(2, 0, 0) AND_115 (c1908_wire_316, {c1908_wire_197_3, c1908_wire_193_2});
nor_n #(2, 0, 0) NOR_32 (c1908_wire_317, {c1908_wire_96_15, c1908_wire_291_5});
and_n #(3, 0, 0) AND_116 (c1908_wire_318, {c1908_wire_319, c1908_wire_311, c1908_wire_216_2});
and_n #(2, 0, 0) AND_117 (c1908_wire_320, {c1908_wire_318_0, c1908_wire_143_1});
and_n #(2, 0, 0) AND_118 (c1908_wire_321, {c1908_wire_318_1, c1908_wire_143_2});
notg #(0, 0) NOT_47 (c1908_wire_319, c1908_wire_96_16);
bufg #(0, 0) BUF_11 (G1884_net_0, c1908_wire_322);
or_n #(2, 0, 0) OR_37 (c1908_wire_322, {c1908_wire_257, c1908_wire_323});
nor_n #(2, 0, 0) NOR_33 (c1908_wire_323, {c1908_wire_258_6, c1908_wire_1_3});
bufg #(0, 0) BUF_12 (G1885_net_0, c1908_wire_324);
or_n #(2, 0, 0) OR_38 (c1908_wire_324, {c1908_wire_259, c1908_wire_325});
nor_n #(2, 0, 0) NOR_34 (c1908_wire_325, {c1908_wire_258_7, c1908_wire_11_3});
bufg #(0, 0) BUF_13 (G1886_net_0, c1908_wire_326);
or_n #(2, 0, 0) OR_39 (c1908_wire_326, {c1908_wire_260, c1908_wire_327});
nor_n #(2, 0, 0) NOR_35 (c1908_wire_327, {c1908_wire_258_8, c1908_wire_12_3});
bufg #(0, 0) BUF_14 (G1887_net_0, c1908_wire_328);
or_n #(2, 0, 0) OR_40 (c1908_wire_328, {c1908_wire_261, c1908_wire_329});
nor_n #(2, 0, 0) NOR_36 (c1908_wire_329, {c1908_wire_258_9, c1908_wire_239_2});
bufg #(0, 0) BUF_15 (G1888_net_0, c1908_wire_330);
or_n #(2, 0, 0) OR_41 (c1908_wire_330, {c1908_wire_69, c1908_wire_331});
nor_n #(2, 0, 0) NOR_37 (c1908_wire_331, {c1908_wire_70_4, c1908_wire_2_5});
bufg #(0, 0) BUF_16 (G1889_net_0, c1908_wire_332);
or_n #(2, 0, 0) OR_42 (c1908_wire_332, {c1908_wire_251, c1908_wire_333});
nor_n #(2, 0, 0) NOR_38 (c1908_wire_333, {c1908_wire_70_5, c1908_wire_21_7});
bufg #(0, 0) BUF_17 (G1890_net_0, c1908_wire_334);
or_n #(2, 0, 0) OR_43 (c1908_wire_334, {c1908_wire_266, c1908_wire_335});
nor_n #(2, 0, 0) NOR_39 (c1908_wire_335, {c1908_wire_70_6, c1908_wire_22_5});
bufg #(0, 0) BUF_18 (G1891_net_0, c1908_wire_336);
or_n #(2, 0, 0) OR_44 (c1908_wire_336, {c1908_wire_276, c1908_wire_337});
nor_n #(2, 0, 0) NOR_40 (c1908_wire_337, {c1908_wire_277_6, c1908_wire_43_3});
bufg #(0, 0) BUF_19 (G1892_net_0, c1908_wire_338);
or_n #(2, 0, 0) OR_45 (c1908_wire_338, {c1908_wire_280, c1908_wire_339});
nor_n #(2, 0, 0) NOR_41 (c1908_wire_339, {c1908_wire_277_7, c1908_wire_41_3});
bufg #(0, 0) BUF_20 (G1893_net_0, c1908_wire_340);
or_n #(2, 0, 0) OR_46 (c1908_wire_340, {c1908_wire_281, c1908_wire_341});
nor_n #(2, 0, 0) NOR_42 (c1908_wire_341, {c1908_wire_277_8, c1908_wire_42_3});
bufg #(0, 0) BUF_21 (G1894_net_0, c1908_wire_342);
or_n #(2, 0, 0) OR_47 (c1908_wire_342, {c1908_wire_278, c1908_wire_343});
nor_n #(2, 0, 0) NOR_43 (c1908_wire_343, {c1908_wire_277_9, c1908_wire_279_1});
bufg #(0, 0) BUF_22 (G1895_net_0, c1908_wire_344);
or_n #(2, 0, 0) OR_48 (c1908_wire_344, {c1908_wire_286, c1908_wire_345});
nor_n #(2, 0, 0) NOR_44 (c1908_wire_345, {c1908_wire_287_2, c1908_wire_15_5});
bufg #(0, 0) BUF_23 (G1896_net_0, c1908_wire_346);
or_n #(2, 0, 0) OR_49 (c1908_wire_346, {c1908_wire_100, c1908_wire_347});
nor_n #(2, 0, 0) NOR_45 (c1908_wire_347, {c1908_wire_101_5, c1908_wire_31_4});
bufg #(0, 0) BUF_24 (G1897_net_0, c1908_wire_348);
or_n #(2, 0, 0) OR_50 (c1908_wire_348, {c1908_wire_146, c1908_wire_349});
nor_n #(2, 0, 0) NOR_46 (c1908_wire_349, {c1908_wire_101_6, c1908_wire_29_5});
bufg #(0, 0) BUF_25 (G1898_net_0, c1908_wire_350);
or_n #(2, 0, 0) OR_51 (c1908_wire_350, {c1908_wire_214, c1908_wire_351});
nor_n #(2, 0, 0) NOR_47 (c1908_wire_351, {c1908_wire_101_7, c1908_wire_30_4});
bufg #(0, 0) BUF_26 (G1899_net_0, c1908_wire_352);
or_n #(2, 0, 0) OR_52 (c1908_wire_352, {c1908_wire_240, c1908_wire_353});
nor_n #(2, 0, 0) NOR_48 (c1908_wire_353, {c1908_wire_101_8, c1908_wire_67_5});
and_n #(3, 0, 0) AND_119 (c1908_wire_252, {c1908_wire_235_4, c1908_wire_354, c1908_wire_355});
bufg #(0, 0) BUF_27 (c1908_wire_197, G19_net_0);
bufg #(0, 0) BUF_28 (G1900_net_0, c1908_wire_356);
notg #(0, 0) NOT_48 (c1908_wire_356, c1908_wire_357);
and_n #(3, 0, 0) AND_120 (c1908_wire_357, {c1908_wire_358, c1908_wire_359, c1908_wire_245});
or_n #(2, 0, 0) OR_53 (c1908_wire_358, {c1908_wire_360, c1908_wire_292});
notg #(0, 0) NOT_49 (c1908_wire_360, c1908_wire_361_0);
notg #(0, 0) NOT_50 (c1908_wire_359, c1908_wire_54_6);
bufg #(0, 0) BUF_29 (G1901_net_0, c1908_wire_362);
nor_n #(2, 0, 0) NOR_49 (c1908_wire_363, {c1908_wire_121_3, c1908_wire_138});
notg #(0, 0) NOT_51 (c1908_wire_364, c1908_wire_365_0);
and_n #(2, 0, 0) AND_121 (c1908_wire_362, {c1908_wire_364, c1908_wire_366});
or_n #(2, 0, 0) OR_54 (c1908_wire_366, {c1908_wire_126, c1908_wire_363});
bufg #(0, 0) BUF_30 (G1902_net_0, c1908_wire_367);
or_n #(2, 0, 0) OR_55 (c1908_wire_368, {c1908_wire_202, c1908_wire_369});
nor_n #(2, 0, 0) NOR_50 (c1908_wire_369, {c1908_wire_200_3, c1908_wire_203_1});
notg #(0, 0) NOT_52 (c1908_wire_370, c1908_wire_365_1);
and_n #(2, 0, 0) AND_122 (c1908_wire_367, {c1908_wire_370, c1908_wire_368});
bufg #(0, 0) BUF_31 (G1903_net_0, c1908_wire_371);
and_n #(2, 0, 0) AND_123 (c1908_wire_371, {c1908_wire_118, c1908_wire_372});
notg #(0, 0) NOT_53 (c1908_wire_372, c1908_wire_365_2);
bufg #(0, 0) BUF_32 (G1904_net_0, c1908_wire_373);
and_n #(2, 0, 0) AND_124 (c1908_wire_373, {c1908_wire_98, c1908_wire_374});
notg #(0, 0) NOT_54 (c1908_wire_374, c1908_wire_365_3);
bufg #(0, 0) BUF_33 (G1905_net_0, c1908_wire_375);
and_n #(2, 0, 0) AND_125 (c1908_wire_375, {c1908_wire_131, c1908_wire_376});
notg #(0, 0) NOT_55 (c1908_wire_376, c1908_wire_365_4);
bufg #(0, 0) BUF_34 (G1906_net_0, c1908_wire_377);
or_n #(2, 0, 0) OR_56 (c1908_wire_149, {c1908_wire_301, c1908_wire_378});
or_n #(2, 0, 0) OR_57 (c1908_wire_379, {c1908_wire_304, c1908_wire_380});
or_n #(2, 0, 0) OR_58 (c1908_wire_377, {c1908_wire_148, c1908_wire_381});
nor_n #(2, 0, 0) NOR_51 (c1908_wire_381, {c1908_wire_379, c1908_wire_135_1});
nor_n #(2, 0, 0) NOR_52 (c1908_wire_378, {c1908_wire_302_2, c1908_wire_303_2});
nor_n #(2, 0, 0) NOR_53 (c1908_wire_380, {c1908_wire_302_3, c1908_wire_303_3});
bufg #(0, 0) BUF_35 (G1907_net_0, c1908_wire_382);
and_n #(2, 0, 0) AND_126 (c1908_wire_383, {c1908_wire_105, c1908_wire_52_2});
notg #(0, 0) NOT_56 (c1908_wire_384, c1908_wire_110);
and_n #(3, 0, 0) AND_127 (c1908_wire_385, {c1908_wire_293, c1908_wire_386, c1908_wire_387_0});
or_n #(2, 0, 0) OR_59 (c1908_wire_295, {c1908_wire_383, c1908_wire_388});
nor_n #(2, 0, 0) NOR_54 (c1908_wire_389, {c1908_wire_107, c1908_wire_52_3});
and_n #(2, 0, 0) AND_128 (c1908_wire_390, {c1908_wire_108, c1908_wire_54_7});
or_n #(3, 0, 0) OR_60 (c1908_wire_382, {c1908_wire_390, c1908_wire_385, c1908_wire_294});
and_n #(2, 0, 0) AND_129 (c1908_wire_391, {c1908_wire_109, c1908_wire_392});
or_n #(2, 0, 0) OR_61 (c1908_wire_386, {c1908_wire_391, c1908_wire_393});
and_n #(2, 0, 0) AND_130 (c1908_wire_394, {c1908_wire_395, c1908_wire_52_4});
and_n #(2, 0, 0) AND_131 (c1908_wire_393, {c1908_wire_394, c1908_wire_384});
or_n #(2, 0, 0) OR_62 (c1908_wire_396, {c1908_wire_389, c1908_wire_397});
and_n #(2, 0, 0) AND_132 (c1908_wire_388, {c1908_wire_396, c1908_wire_398});
notg #(0, 0) NOT_57 (c1908_wire_397, c1908_wire_387_1);
notg #(0, 0) NOT_58 (c1908_wire_398, c1908_wire_54_8);
notg #(0, 0) NOT_59 (c1908_wire_392, c1908_wire_52_5);
notg #(0, 0) NOT_60 (c1908_wire_395, c1908_wire_54_9);
bufg #(0, 0) BUF_36 (G1908_net_0, c1908_wire_399);
or_n #(2, 0, 0) OR_63 (c1908_wire_145, {c1908_wire_320, c1908_wire_400});
nor_n #(2, 0, 0) NOR_55 (c1908_wire_401, {c1908_wire_318_2, c1908_wire_143_3});
or_n #(2, 0, 0) OR_64 (c1908_wire_402, {c1908_wire_401, c1908_wire_321});
or_n #(2, 0, 0) OR_65 (c1908_wire_403, {c1908_wire_144, c1908_wire_404});
nor_n #(2, 0, 0) NOR_56 (c1908_wire_404, {c1908_wire_402, c1908_wire_140_2});
and_n #(2, 0, 0) AND_133 (c1908_wire_399, {c1908_wire_403, c1908_wire_405});
nor_n #(2, 0, 0) NOR_57 (c1908_wire_400, {c1908_wire_318_3, c1908_wire_143_4});
notg #(0, 0) NOT_61 (c1908_wire_405, c1908_wire_365_5);
and_n #(3, 0, 0) AND_134 (c1908_wire_79, {c1908_wire_197_4, c1908_wire_406, c1908_wire_407});
xor_n #(2, 0, 0) XOR_35 (c1908_wire_143, {c1908_wire_1_4, c1908_wire_296});
bufg #(0, 0) BUF_37 (c1908_wire_11, G2_net_0);
bufg #(0, 0) BUF_38 (c1908_wire_408, G20_net_0);
and_n #(2, 0, 0) AND_135 (c1908_wire_169, {c1908_wire_408_0, c1908_wire_409});
and_n #(3, 0, 0) AND_136 (c1908_wire_213, {c1908_wire_408_1, c1908_wire_410, c1908_wire_411});
bufg #(0, 0) BUF_39 (c1908_wire_85, G21_net_0);
bufg #(0, 0) BUF_40 (c1908_wire_52, G22_net_0);
bufg #(0, 0) BUF_41 (c1908_wire_193, G23_net_0);
notg #(0, 0) NOT_62 (c1908_wire_412, c1908_wire_193_3);
notg #(0, 0) NOT_63 (c1908_wire_406, c1908_wire_193_4);
notg #(0, 0) NOT_64 (c1908_wire_410, c1908_wire_193_5);
bufg #(0, 0) BUF_42 (c1908_wire_300, G24_net_0);
and_n #(2, 0, 0) AND_137 (c1908_wire_413, {c1908_wire_300_1, c1908_wire_412});
notg #(0, 0) NOT_65 (c1908_wire_297, c1908_wire_300_2);
notg #(0, 0) NOT_66 (c1908_wire_354, c1908_wire_300_3);
bufg #(0, 0) BUF_43 (c1908_wire_231, G25_net_0);
bufg #(0, 0) BUF_44 (c1908_wire_216, G26_net_0);
bufg #(0, 0) BUF_45 (c1908_wire_183, G27_net_0);
bufg #(0, 0) BUF_46 (c1908_wire_172, G28_net_0);
bufg #(0, 0) BUF_47 (c1908_wire_150, G29_net_0);
and_n #(2, 0, 0) AND_138 (c1908_wire_414, {c1908_wire_11_4, c1908_wire_415});
bufg #(0, 0) BUF_48 (c1908_wire_12, G3_net_0);
bufg #(0, 0) BUF_49 (c1908_wire_387, G30_net_0);
bufg #(0, 0) BUF_50 (c1908_wire_96, G31_net_0);
bufg #(0, 0) BUF_51 (c1908_wire_361, G32_net_0);
nor_n #(2, 0, 0) NOR_58 (c1908_wire_365, {c1908_wire_361_1, c1908_wire_54_10});
bufg #(0, 0) BUF_52 (c1908_wire_54, G33_net_0);
notg #(0, 0) NOT_67 (c1908_wire_298, c1908_wire_54_11);
notg #(0, 0) NOT_68 (c1908_wire_407, c1908_wire_54_12);
notg #(0, 0) NOT_69 (c1908_wire_411, c1908_wire_54_13);
notg #(0, 0) NOT_70 (c1908_wire_355, c1908_wire_54_14);
notg #(0, 0) NOT_71 (c1908_wire_416, c1908_wire_54_15);
nor_n #(2, 0, 0) NOR_59 (c1908_wire_417, {c1908_wire_193_6, c1908_wire_96_17});
notg #(0, 0) NOT_72 (c1908_wire_409, c1908_wire_417);
nor_n #(2, 0, 0) NOR_60 (c1908_wire_237, {c1908_wire_300_4, c1908_wire_96_18});
and_n #(2, 0, 0) AND_139 (c1908_wire_418, {c1908_wire_12_4, c1908_wire_419});
bufg #(0, 0) BUF_53 (c1908_wire_239, G4_net_0);
and_n #(2, 0, 0) AND_140 (c1908_wire_303, {c1908_wire_416, c1908_wire_420});
nand_n #(2, 0, 0) NAND_1 (c1908_wire_420, {c1908_wire_85_2, c1908_wire_150_1});
and_n #(2, 0, 0) AND_141 (c1908_wire_421, {c1908_wire_239_3, c1908_wire_279_2});
xor_n #(2, 0, 0) XOR_36 (c1908_wire_72, {c1908_wire_239_4, c1908_wire_42_4});
xor_n #(2, 0, 0) XOR_37 (c1908_wire_422, {c1908_wire_239_5, c1908_wire_42_5});
bufg #(0, 0) BUF_54 (c1908_wire_43, G5_net_0);
nor_n #(4, 0, 0) NOR_61 (c1908_wire_423, {c1908_wire_150_2, c1908_wire_96_19, c1908_wire_54_16, c1908_wire_413_0});
nor_n #(4, 0, 0) NOR_62 (c1908_wire_424, {c1908_wire_387_2, c1908_wire_96_20, c1908_wire_54_17, c1908_wire_413_1});
nor_n #(3, 0, 0) NOR_63 (c1908_wire_163, {c1908_wire_54_18, c1908_wire_361_2, c1908_wire_413_2});
xor_n #(2, 0, 0) XOR_38 (c1908_wire_415, {c1908_wire_43_4, c1908_wire_279_3});
xor_n #(2, 0, 0) XOR_39 (c1908_wire_425, {c1908_wire_43_5, c1908_wire_279_4});
bufg #(0, 0) BUF_55 (c1908_wire_41, G6_net_0);
xor_n #(2, 0, 0) XOR_40 (c1908_wire_419, {c1908_wire_41_4, c1908_wire_279_5});
xor_n #(2, 0, 0) XOR_41 (c1908_wire_426, {c1908_wire_41_5, c1908_wire_279_6});
bufg #(0, 0) BUF_56 (c1908_wire_42, G7_net_0);
or_n #(2, 0, 0) OR_66 (c1908_wire_36, {c1908_wire_421, c1908_wire_427});
nor_n #(2, 0, 0) NOR_64 (c1908_wire_427, {c1908_wire_279_7, c1908_wire_239_6});
or_n #(2, 0, 0) OR_67 (c1908_wire_106, {c1908_wire_238, c1908_wire_428});
nor_n #(2, 0, 0) NOR_65 (c1908_wire_428, {c1908_wire_67_6, c1908_wire_15_6});
or_n #(2, 0, 0) OR_68 (c1908_wire_111, {c1908_wire_212, c1908_wire_429});
nor_n #(2, 0, 0) NOR_66 (c1908_wire_429, {c1908_wire_213_1, c1908_wire_30_5});
nor_n #(2, 0, 0) NOR_67 (c1908_wire_265, {c1908_wire_423, c1908_wire_163_3});
nor_n #(2, 0, 0) NOR_68 (c1908_wire_268, {c1908_wire_424, c1908_wire_163_4});
bufg #(0, 0) BUF_57 (c1908_wire_279, G8_net_0);
bufg #(0, 0) BUF_58 (c1908_wire_15, G9_net_0);
nor_n #(2, 0, 0) NOR_69 (c1908_wire_430, {c1908_wire_2_6, c1908_wire_422});
or_n #(2, 0, 0) OR_69 (c1908_wire_112, {c1908_wire_71, c1908_wire_430});
nor_n #(2, 0, 0) NOR_70 (c1908_wire_431, {c1908_wire_11_5, c1908_wire_425});
or_n #(2, 0, 0) OR_70 (c1908_wire_87, {c1908_wire_414, c1908_wire_431});
nor_n #(2, 0, 0) NOR_71 (c1908_wire_432, {c1908_wire_31_5, c1908_wire_253});
or_n #(2, 0, 0) OR_71 (c1908_wire_88, {c1908_wire_102, c1908_wire_432});
nor_n #(2, 0, 0) NOR_72 (c1908_wire_433, {c1908_wire_2_7, c1908_wire_147});
or_n #(2, 0, 0) OR_72 (c1908_wire_76, {c1908_wire_73, c1908_wire_433});
nor_n #(2, 0, 0) NOR_73 (c1908_wire_434, {c1908_wire_12_5, c1908_wire_426});
or_n #(2, 0, 0) OR_73 (c1908_wire_77, {c1908_wire_418, c1908_wire_434});

endmodule
