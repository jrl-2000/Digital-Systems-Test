// Fanout-inserted! -- Created by V2S
// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module c1908_fo (N1_PI,N4_PI,N7_PI,N10_PI,N13_PI,N16_PI,N19_PI,N22_PI,N25_PI,N28_PI,
              N31_PI,N34_PI,N37_PI,N40_PI,N43_PI,N46_PI,N49_PI,N53_PI,N56_PI,N60_PI,
              N63_PI,N66_PI,N69_PI,N72_PI,N76_PI,N79_PI,N82_PI,N85_PI,N88_PI,N91_PI,
              N94_PI,N99_PI,N104_PI,N2753_PO,N2754_PO,N2755_PO,N2756_PO,N2762_PO,N2767_PO,N2768_PO,
              N2779_PO,N2780_PO,N2781_PO,N2782_PO,N2783_PO,N2784_PO,N2785_PO,N2786_PO,N2787_PO,N2811_PO,
              N2886_PO,N2887_PO,N2888_PO,N2889_PO,N2890_PO,N2891_PO,N2892_PO,N2899_PO);

input N1_PI,N4_PI,N7_PI,N10_PI,N13_PI,N16_PI,N19_PI,N22_PI,N25_PI,N28_PI,
      N31_PI,N34_PI,N37_PI,N40_PI,N43_PI,N46_PI,N49_PI,N53_PI,N56_PI,N60_PI,
      N63_PI,N66_PI,N69_PI,N72_PI,N76_PI,N79_PI,N82_PI,N85_PI,N88_PI,N91_PI,
      N94_PI,N99_PI,N104_PI;

output N2753_PO,N2754_PO,N2755_PO,N2756_PO,N2762_PO,N2767_PO,N2768_PO,N2779_PO,N2780_PO,N2781_PO,
       N2782_PO,N2783_PO,N2784_PO,N2785_PO,N2786_PO,N2787_PO,N2811_PO,N2886_PO,N2887_PO,N2888_PO,
       N2889_PO,N2890_PO,N2891_PO,N2892_PO,N2899_PO;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898;

// New Introduced Signals (inputs/outputs)
wire N1, N4, N7, N10, N13, N16, N19, 
     N22, N25, N28, N31, N34, N37, N40, N43, 
     N46, N49, N53, N56, N60, N63, N66, N69, 
     N72, N76, N79, N82, N85, N88, N91, N94, 
     N99, N104, N2753, N2754, N2755, N2756, N2762, N2767, 
     N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, 
     N2786, N2787, N2811, N2886, N2887, N2888, N2889, N2890, 
     N2891, N2892, N2899;

// New Introduced Signals (fanouts)
wire N1_0, N1_1,
     N4_0, N4_1,
     N7_0, N7_1,
     N10_0, N10_1,
     N13_0, N13_1,
     N16_0, N16_1,
     N19_0, N19_1,
     N22_0, N22_1,
     N25_0, N25_1,
     N28_0, N28_1,
     N31_0, N31_1,
     N34_0, N34_1,
     N37_0, N37_1,
     N40_0, N40_1,
     N43_0, N43_1,
     N46_0, N46_1,
     N49_0, N49_1, N49_2,
     N53_0, N53_1,
     N56_0, N56_1, N56_2,
     N60_0, N60_1,
     N63_0, N63_1,
     N66_0, N66_1,
     N69_0, N69_1,
     N72_0, N72_1, N72_2,
     N76_0, N76_1,
     N79_0, N79_1,
     N82_0, N82_1,
     N85_0, N85_1,
     N88_0, N88_1,
     N91_0, N91_1,
     N94_0, N94_1, N94_2, N94_3,
     N99_0, N99_1, N99_2, N99_3,
     N104_0, N104_1, N104_2, N104_3, N104_4, N104_5, N104_6,
     N190_0, N190_1, N190_2,
     N194_0, N194_1,
     N197_0, N197_1, N197_2,
     N201_0, N201_1, N201_2, N201_3,
     N206_0, N206_1,
     N209_0, N209_1,
     N212_0, N212_1, N212_2,
     N216_0, N216_1, N216_2,
     N220_0, N220_1, N220_2, N220_3,
     N225_0, N225_1, N225_2,
     N229_0, N229_1,
     N232_0, N232_1,
     N235_0, N235_1, N235_2,
     N239_0, N239_1, N239_2,
     N243_0, N243_1, N243_2,
     N247_0, N247_1, N247_2,
     N253_0, N253_1,
     N257_0, N257_1,
     N260_0, N260_1,
     N263_0, N263_1,
     N266_0, N266_1,
     N269_0, N269_1,
     N272_0, N272_1,
     N277_0, N277_1,
     N280_0, N280_1,
     N283_0, N283_1, N283_2, N283_3, N283_4, N283_5,
     N290_0, N290_1, N290_2, N290_3, N290_4, N290_5,
     N297_0, N297_1,
     N300_0, N300_1,
     N303_0, N303_1,
     N306_0, N306_1, N306_2, N306_3, N306_4, N306_5,
     N313_0, N313_1,
     N316_0, N316_1,
     N319_0, N319_1, N319_2, N319_3, N319_4, N319_5,
     N326_0, N326_1, N326_2, N326_3,
     N331_0, N331_1, N331_2, N331_3, N331_4, N331_5,
     N338_0, N338_1, N338_2, N338_3,
     N343_0, N343_1,
     N346_0, N346_1,
     N349_0, N349_1,
     N352_0, N352_1,
     N355_0, N355_1,
     N358_0, N358_1,
     N361_0, N361_1,
     N364_0, N364_1,
     N367_0, N367_1,
     N370_0, N370_1,
     N373_0, N373_1,
     N376_0, N376_1,
     N379_0, N379_1,
     N382_0, N382_1,
     N385_0, N385_1,
     N388_0, N388_1,
     N556_0, N556_1,
     N559_0, N559_1,
     N562_0, N562_1,
     N565_0, N565_1,
     N568_0, N568_1,
     N571_0, N571_1,
     N574_0, N574_1,
     N577_0, N577_1,
     N580_0, N580_1,
     N583_0, N583_1,
     N586_0, N586_1,
     N589_0, N589_1,
     N592_0, N592_1,
     N595_0, N595_1,
     N598_0, N598_1,
     N603_0, N603_1, N603_2, N603_3,
     N608_0, N608_1, N608_2,
     N612_0, N612_1, N612_2,
     N616_0, N616_1,
     N619_0, N619_1,
     N622_0, N622_1,
     N625_0, N625_1,
     N628_0, N628_1,
     N631_0, N631_1,
     N634_0, N634_1,
     N637_0, N637_1,
     N640_0, N640_1,
     N643_0, N643_1,
     N646_0, N646_1,
     N649_0, N649_1,
     N652_0, N652_1,
     N655_0, N655_1,
     N658_0, N658_1,
     N661_0, N661_1,
     N664_0, N664_1,
     N667_0, N667_1,
     N670_0, N670_1,
     N673_0, N673_1,
     N676_0, N676_1,
     N679_0, N679_1,
     N682_0, N682_1,
     N685_0, N685_1,
     N688_0, N688_1,
     N691_0, N691_1,
     N694_0, N694_1,
     N697_0, N697_1,
     N700_0, N700_1,
     N703_0, N703_1,
     N706_0, N706_1,
     N709_0, N709_1,
     N712_0, N712_1,
     N715_0, N715_1,
     N718_0, N718_1,
     N721_0, N721_1,
     N724_0, N724_1,
     N727_0, N727_1,
     N730_0, N730_1,
     N733_0, N733_1,
     N736_0, N736_1,
     N739_0, N739_1,
     N742_0, N742_1,
     N745_0, N745_1,
     N748_0, N748_1,
     N751_0, N751_1,
     N899_0, N899_1, N899_2,
     N903_0, N903_1, N903_2,
     N907_0, N907_1,
     N910_0, N910_1,
     N923_0, N923_1,
     N926_0, N926_1, N926_2, N926_3, N926_4, N926_5, N926_6, N926_7,
     N935_0, N935_1,
     N939_0, N939_1,
     N943_0, N943_1,
     N947_0, N947_1,
     N951_0, N951_1,
     N955_0, N955_1,
     N959_0, N959_1,
     N962_0, N962_1,
     N965_0, N965_1,
     N969_0, N969_1,
     N973_0, N973_1,
     N977_0, N977_1,
     N981_0, N981_1,
     N985_0, N985_1,
     N994_0, N994_1,
     N998_0, N998_1,
     N1010_0, N1010_1,
     N1013_0, N1013_1,
     N1016_0, N1016_1,
     N1019_0, N1019_1,
     N1022_0, N1022_1,
     N1025_0, N1025_1,
     N1028_0, N1028_1,
     N1031_0, N1031_1,
     N1034_0, N1034_1,
     N1037_0, N1037_1,
     N1040_0, N1040_1,
     N1043_0, N1043_1,
     N1046_0, N1046_1,
     N1049_0, N1049_1,
     N1164_0, N1164_1,
     N1168_0, N1168_1,
     N1171_0, N1171_1, N1171_2, N1171_3, N1171_4, N1171_5, N1171_6, N1171_7, N1171_8, N1171_9, N1171_10, N1171_11, N1171_12, N1171_13, N1171_14, N1171_15,
     N1188_0, N1188_1, N1188_2, N1188_3, N1188_4, N1188_5, N1188_6, N1188_7, N1188_8, N1188_9, N1188_10, N1188_11, N1188_12, N1188_13, N1188_14, N1188_15,
     N1232_0, N1232_1,
     N1235_0, N1235_1,
     N1243_0, N1243_1,
     N1246_0, N1246_1,
     N1249_0, N1249_1,
     N1252_0, N1252_1,
     N1255_0, N1255_1,
     N1258_0, N1258_1,
     N1261_0, N1261_1,
     N1264_0, N1264_1,
     N1319_0, N1319_1,
     N1334_0, N1334_1,
     N1352_0, N1352_1,
     N1355_0, N1355_1,
     N1358_0, N1358_1,
     N1361_0, N1361_1,
     N1364_0, N1364_1,
     N1367_0, N1367_1,
     N1370_0, N1370_1,
     N1373_0, N1373_1,
     N1376_0, N1376_1,
     N1379_0, N1379_1,
     N1383_0, N1383_1,
     N1390_0, N1390_1,
     N1393_0, N1393_1,
     N1416_0, N1416_1,
     N1419_0, N1419_1,
     N1440_0, N1440_1,
     N1472_0, N1472_1,
     N1478_0, N1478_1,
     N1481_0, N1481_1,
     N1484_0, N1484_1,
     N1510_0, N1510_1,
     N1514_0, N1514_1,
     N1517_0, N1517_1,
     N1522_0, N1522_1, N1522_2,
     N1534_0, N1534_1,
     N1537_0, N1537_1,
     N1540_0, N1540_1,
     N1546_0, N1546_1,
     N1554_0, N1554_1,
     N1557_0, N1557_1, N1557_2,
     N1561_0, N1561_1,
     N1571_0, N1571_1,
     N1576_0, N1576_1,
     N1588_0, N1588_1,
     N1596_0, N1596_1,
     N1600_0, N1600_1,
     N1603_0, N1603_1,
     N1606_0, N1606_1,
     N1609_0, N1609_1,
     N1612_0, N1612_1,
     N1615_0, N1615_1,
     N1620_0, N1620_1,
     N1623_0, N1623_1,
     N1640_0, N1640_1,
     N1643_0, N1643_1,
     N1647_0, N1647_1,
     N1651_0, N1651_1,
     N1658_0, N1658_1,
     N1661_0, N1661_1,
     N1664_0, N1664_1,
     N1685_0, N1685_1,
     N1697_0, N1697_1,
     N1701_0, N1701_1,
     N1714_0, N1714_1,
     N1717_0, N1717_1,
     N1723_0, N1723_1,
     N1731_0, N1731_1,
     N1734_0, N1734_1,
     N1742_0, N1742_1,
     N1748_0, N1748_1,
     N1751_0, N1751_1,
     N1774_0, N1774_1,
     N1777_0, N1777_1,
     N1788_0, N1788_1,
     N1798_0, N1798_1,
     N1802_0, N1802_1,
     N1812_0, N1812_1,
     N1815_0, N1815_1,
     N1818_0, N1818_1,
     N1830_0, N1830_1,
     N1838_0, N1838_1,
     N1841_0, N1841_1,
     N1858_0, N1858_1,
     N1866_0, N1866_1,
     N1869_0, N1869_1,
     N1872_0, N1872_1,
     N1875_0, N1875_1,
     N1879_0, N1879_1,
     N1889_0, N1889_1,
     N1898_0, N1898_1,
     N1902_0, N1902_1,
     N1927_0, N1927_1,
     N1930_0, N1930_1,
     N1933_0, N1933_1,
     N1944_0, N1944_1,
     N1947_0, N1947_1,
     N1950_0, N1950_1,
     N1953_0, N1953_1,
     N1958_0, N1958_1,
     N1961_0, N1961_1,
     N1965_0, N1965_1,
     N1968_0, N1968_1,
     N1980_0, N1980_1,
     N1987_0, N1987_1,
     N2027_0, N2027_1,
     N2030_0, N2030_1,
     N2033_0, N2033_1,
     N2042_0, N2042_1,
     N2052_0, N2052_1,
     N2055_0, N2055_1,
     N2062_0, N2062_1,
     N2068_0, N2068_1,
     N2071_0, N2071_1,
     N2078_0, N2078_1,
     N2081_0, N2081_1,
     N2086_0, N2086_1,
     N2089_0, N2089_1,
     N2104_0, N2104_1, N2104_2, N2104_3, N2104_4, N2104_5, N2104_6, N2104_7, N2104_8, N2104_9, N2104_10, N2104_11, N2104_12, N2104_13,
     N2119_0, N2119_1, N2119_2, N2119_3, N2119_4, N2119_5, N2119_6, N2119_7, N2119_8,
     N2129_0, N2129_1, N2129_2, N2129_3, N2129_4, N2129_5, N2129_6, N2129_7, N2129_8, N2129_9, N2129_10, N2129_11, N2129_12,
     N2143_0, N2143_1, N2143_2, N2143_3,
     N2148_0, N2148_1,
     N2151_0, N2151_1,
     N2196_0, N2196_1,
     N2199_0, N2199_1,
     N2202_0, N2202_1,
     N2205_0, N2205_1,
     N2237_0, N2237_1,
     N2241_0, N2241_1,
     N2245_0, N2245_1,
     N2257_0, N2257_1,
     N2260_0, N2260_1,
     N2263_0, N2263_1,
     N2266_0, N2266_1,
     N2269_0, N2269_1,
     N2272_0, N2272_1,
     N2279_0, N2279_1,
     N2286_0, N2286_1, N2286_2, N2286_3, N2286_4, N2286_5, N2286_6, N2286_7, N2286_8, N2286_9,
     N2297_0, N2297_1, N2297_2, N2297_3, N2297_4, N2297_5, N2297_6, N2297_7, N2297_8, N2297_9, N2297_10, N2297_11, N2297_12, N2297_13, N2297_14,
     N2315_0, N2315_1, N2315_2, N2315_3, N2315_4, N2315_5, N2315_6, N2315_7, N2315_8, N2315_9,
     N2326_0, N2326_1, N2326_2, N2326_3, N2326_4, N2326_5, N2326_6, N2326_7, N2326_8, N2326_9, N2326_10, N2326_11, N2326_12,
     N2340_0, N2340_1, N2340_2, N2340_3, N2340_4, N2340_5, N2340_6, N2340_7, N2340_8, N2340_9, N2340_10, N2340_11,
     N2353_0, N2353_1, N2353_2, N2353_3, N2353_4, N2353_5, N2353_6,
     N2361_0, N2361_1, N2361_2, N2361_3, N2361_4, N2361_5, N2361_6, N2361_7, N2361_8, N2361_9, N2361_10, N2361_11, N2361_12,
     N2375_0, N2375_1, N2375_2, N2375_3, N2375_4, N2375_5, N2375_6, N2375_7,
     N2386_0, N2386_1, N2386_2, N2386_3, N2386_4, N2386_5, N2386_6, N2386_7, N2386_8, N2386_9, N2386_10, N2386_11, N2386_12, N2386_13,
     N2427_0, N2427_1, N2427_2, N2427_3, N2427_4, N2427_5, N2427_6, N2427_7, N2427_8, N2427_9, N2427_10, N2427_11, N2427_12, N2427_13, N2427_14, N2427_15,
     N2537_0, N2537_1,
     N2540_0, N2540_1,
     N2543_0, N2543_1,
     N2546_0, N2546_1,
     N2549_0, N2549_1,
     N2552_0, N2552_1,
     N2555_0, N2555_1,
     N2558_0, N2558_1,
     N2561_0, N2561_1,
     N2564_0, N2564_1,
     N2567_0, N2567_1,
     N2570_0, N2570_1,
     N2573_0, N2573_1,
     N2576_0, N2576_1,
     N2594_0, N2594_1,
     N2597_0, N2597_1,
     N2600_0, N2600_1,
     N2603_0, N2603_1,
     N2606_0, N2606_1,
     N2611_0, N2611_1,
     N2614_0, N2614_1,
     N2617_0, N2617_1,
     N2620_0, N2620_1,
     N2639_0, N2639_1,
     N2642_0, N2642_1,
     N2645_0, N2645_1,
     N2648_0, N2648_1,
     N2651_0, N2651_1,
     N2655_0, N2655_1,
     N2658_0, N2658_1,
     N2661_0, N2661_1,
     N2664_0, N2664_1,
     N2747_0, N2747_1,
     N2750_0, N2750_1,
     N2773_0, N2773_1,
     N2776_0, N2776_1,
     N2789_0, N2789_1, N2789_2, N2789_3, N2789_4, N2789_5,
     N2812_0, N2812_1,
     N2815_0, N2815_1,
     N2818_0, N2818_1,
     N2821_0, N2821_1,
     N2824_0, N2824_1,
     N2829_0, N2829_1,
     N2843_0, N2843_1,
     N2846_0, N2846_1,
     N2883_0, N2883_1;

// New Primary Input (PI) components
pin pin_0 (N1_PI, N1);
pin pin_1 (N4_PI, N4);
pin pin_2 (N7_PI, N7);
pin pin_3 (N10_PI, N10);
pin pin_4 (N13_PI, N13);
pin pin_5 (N16_PI, N16);
pin pin_6 (N19_PI, N19);
pin pin_7 (N22_PI, N22);
pin pin_8 (N25_PI, N25);
pin pin_9 (N28_PI, N28);
pin pin_10 (N31_PI, N31);
pin pin_11 (N34_PI, N34);
pin pin_12 (N37_PI, N37);
pin pin_13 (N40_PI, N40);
pin pin_14 (N43_PI, N43);
pin pin_15 (N46_PI, N46);
pin pin_16 (N49_PI, N49);
pin pin_17 (N53_PI, N53);
pin pin_18 (N56_PI, N56);
pin pin_19 (N60_PI, N60);
pin pin_20 (N63_PI, N63);
pin pin_21 (N66_PI, N66);
pin pin_22 (N69_PI, N69);
pin pin_23 (N72_PI, N72);
pin pin_24 (N76_PI, N76);
pin pin_25 (N79_PI, N79);
pin pin_26 (N82_PI, N82);
pin pin_27 (N85_PI, N85);
pin pin_28 (N88_PI, N88);
pin pin_29 (N91_PI, N91);
pin pin_30 (N94_PI, N94);
pin pin_31 (N99_PI, N99);
pin pin_32 (N104_PI, N104);

// New Primary Output (PO) components
pout pout_0 (N2753, N2753_PO);
pout pout_1 (N2754, N2754_PO);
pout pout_2 (N2755, N2755_PO);
pout pout_3 (N2756, N2756_PO);
pout pout_4 (N2762, N2762_PO);
pout pout_5 (N2767, N2767_PO);
pout pout_6 (N2768, N2768_PO);
pout pout_7 (N2779, N2779_PO);
pout pout_8 (N2780, N2780_PO);
pout pout_9 (N2781, N2781_PO);
pout pout_10 (N2782, N2782_PO);
pout pout_11 (N2783, N2783_PO);
pout pout_12 (N2784, N2784_PO);
pout pout_13 (N2785, N2785_PO);
pout pout_14 (N2786, N2786_PO);
pout pout_15 (N2787, N2787_PO);
pout pout_16 (N2811, N2811_PO);
pout pout_17 (N2886, N2886_PO);
pout pout_18 (N2887, N2887_PO);
pout pout_19 (N2888, N2888_PO);
pout pout_20 (N2889, N2889_PO);
pout pout_21 (N2890, N2890_PO);
pout pout_22 (N2891, N2891_PO);
pout pout_23 (N2892, N2892_PO);
pout pout_24 (N2899, N2899_PO);

// New Fan-out (FANOUT) components
fanout_n #(2,0,0) fanout_n_0 (N1, {N1_0, N1_1});
fanout_n #(2,0,0) fanout_n_1 (N4, {N4_0, N4_1});
fanout_n #(2,0,0) fanout_n_2 (N7, {N7_0, N7_1});
fanout_n #(2,0,0) fanout_n_3 (N10, {N10_0, N10_1});
fanout_n #(2,0,0) fanout_n_4 (N13, {N13_0, N13_1});
fanout_n #(2,0,0) fanout_n_5 (N16, {N16_0, N16_1});
fanout_n #(2,0,0) fanout_n_6 (N19, {N19_0, N19_1});
fanout_n #(2,0,0) fanout_n_7 (N22, {N22_0, N22_1});
fanout_n #(2,0,0) fanout_n_8 (N25, {N25_0, N25_1});
fanout_n #(2,0,0) fanout_n_9 (N28, {N28_0, N28_1});
fanout_n #(2,0,0) fanout_n_10 (N31, {N31_0, N31_1});
fanout_n #(2,0,0) fanout_n_11 (N34, {N34_0, N34_1});
fanout_n #(2,0,0) fanout_n_12 (N37, {N37_0, N37_1});
fanout_n #(2,0,0) fanout_n_13 (N40, {N40_0, N40_1});
fanout_n #(2,0,0) fanout_n_14 (N43, {N43_0, N43_1});
fanout_n #(2,0,0) fanout_n_15 (N46, {N46_0, N46_1});
fanout_n #(3,0,0) fanout_n_16 (N49, {N49_0, N49_1, N49_2});
fanout_n #(2,0,0) fanout_n_17 (N53, {N53_0, N53_1});
fanout_n #(3,0,0) fanout_n_18 (N56, {N56_0, N56_1, N56_2});
fanout_n #(2,0,0) fanout_n_19 (N60, {N60_0, N60_1});
fanout_n #(2,0,0) fanout_n_20 (N63, {N63_0, N63_1});
fanout_n #(2,0,0) fanout_n_21 (N66, {N66_0, N66_1});
fanout_n #(2,0,0) fanout_n_22 (N69, {N69_0, N69_1});
fanout_n #(3,0,0) fanout_n_23 (N72, {N72_0, N72_1, N72_2});
fanout_n #(2,0,0) fanout_n_24 (N76, {N76_0, N76_1});
fanout_n #(2,0,0) fanout_n_25 (N79, {N79_0, N79_1});
fanout_n #(2,0,0) fanout_n_26 (N82, {N82_0, N82_1});
fanout_n #(2,0,0) fanout_n_27 (N85, {N85_0, N85_1});
fanout_n #(2,0,0) fanout_n_28 (N88, {N88_0, N88_1});
fanout_n #(2,0,0) fanout_n_29 (N91, {N91_0, N91_1});
fanout_n #(4,0,0) fanout_n_30 (N94, {N94_0, N94_1, N94_2, N94_3});
fanout_n #(4,0,0) fanout_n_31 (N99, {N99_0, N99_1, N99_2, N99_3});
fanout_n #(7,0,0) fanout_n_32 (N104, {N104_0, N104_1, N104_2, N104_3, N104_4, N104_5, N104_6});
fanout_n #(3,0,0) fanout_n_33 (N190, {N190_0, N190_1, N190_2});
fanout_n #(2,0,0) fanout_n_34 (N194, {N194_0, N194_1});
fanout_n #(3,0,0) fanout_n_35 (N197, {N197_0, N197_1, N197_2});
fanout_n #(4,0,0) fanout_n_36 (N201, {N201_0, N201_1, N201_2, N201_3});
fanout_n #(2,0,0) fanout_n_37 (N206, {N206_0, N206_1});
fanout_n #(2,0,0) fanout_n_38 (N209, {N209_0, N209_1});
fanout_n #(3,0,0) fanout_n_39 (N212, {N212_0, N212_1, N212_2});
fanout_n #(3,0,0) fanout_n_40 (N216, {N216_0, N216_1, N216_2});
fanout_n #(4,0,0) fanout_n_41 (N220, {N220_0, N220_1, N220_2, N220_3});
fanout_n #(3,0,0) fanout_n_42 (N225, {N225_0, N225_1, N225_2});
fanout_n #(2,0,0) fanout_n_43 (N229, {N229_0, N229_1});
fanout_n #(2,0,0) fanout_n_44 (N232, {N232_0, N232_1});
fanout_n #(3,0,0) fanout_n_45 (N235, {N235_0, N235_1, N235_2});
fanout_n #(3,0,0) fanout_n_46 (N239, {N239_0, N239_1, N239_2});
fanout_n #(3,0,0) fanout_n_47 (N243, {N243_0, N243_1, N243_2});
fanout_n #(3,0,0) fanout_n_48 (N247, {N247_0, N247_1, N247_2});
fanout_n #(2,0,0) fanout_n_49 (N253, {N253_0, N253_1});
fanout_n #(2,0,0) fanout_n_50 (N257, {N257_0, N257_1});
fanout_n #(2,0,0) fanout_n_51 (N260, {N260_0, N260_1});
fanout_n #(2,0,0) fanout_n_52 (N263, {N263_0, N263_1});
fanout_n #(2,0,0) fanout_n_53 (N266, {N266_0, N266_1});
fanout_n #(2,0,0) fanout_n_54 (N269, {N269_0, N269_1});
fanout_n #(2,0,0) fanout_n_55 (N272, {N272_0, N272_1});
fanout_n #(2,0,0) fanout_n_56 (N277, {N277_0, N277_1});
fanout_n #(2,0,0) fanout_n_57 (N280, {N280_0, N280_1});
fanout_n #(6,0,0) fanout_n_58 (N283, {N283_0, N283_1, N283_2, N283_3, N283_4, N283_5});
fanout_n #(6,0,0) fanout_n_59 (N290, {N290_0, N290_1, N290_2, N290_3, N290_4, N290_5});
fanout_n #(2,0,0) fanout_n_60 (N297, {N297_0, N297_1});
fanout_n #(2,0,0) fanout_n_61 (N300, {N300_0, N300_1});
fanout_n #(2,0,0) fanout_n_62 (N303, {N303_0, N303_1});
fanout_n #(6,0,0) fanout_n_63 (N306, {N306_0, N306_1, N306_2, N306_3, N306_4, N306_5});
fanout_n #(2,0,0) fanout_n_64 (N313, {N313_0, N313_1});
fanout_n #(2,0,0) fanout_n_65 (N316, {N316_0, N316_1});
fanout_n #(6,0,0) fanout_n_66 (N319, {N319_0, N319_1, N319_2, N319_3, N319_4, N319_5});
fanout_n #(4,0,0) fanout_n_67 (N326, {N326_0, N326_1, N326_2, N326_3});
fanout_n #(6,0,0) fanout_n_68 (N331, {N331_0, N331_1, N331_2, N331_3, N331_4, N331_5});
fanout_n #(4,0,0) fanout_n_69 (N338, {N338_0, N338_1, N338_2, N338_3});
fanout_n #(2,0,0) fanout_n_70 (N343, {N343_0, N343_1});
fanout_n #(2,0,0) fanout_n_71 (N346, {N346_0, N346_1});
fanout_n #(2,0,0) fanout_n_72 (N349, {N349_0, N349_1});
fanout_n #(2,0,0) fanout_n_73 (N352, {N352_0, N352_1});
fanout_n #(2,0,0) fanout_n_74 (N355, {N355_0, N355_1});
fanout_n #(2,0,0) fanout_n_75 (N358, {N358_0, N358_1});
fanout_n #(2,0,0) fanout_n_76 (N361, {N361_0, N361_1});
fanout_n #(2,0,0) fanout_n_77 (N364, {N364_0, N364_1});
fanout_n #(2,0,0) fanout_n_78 (N367, {N367_0, N367_1});
fanout_n #(2,0,0) fanout_n_79 (N370, {N370_0, N370_1});
fanout_n #(2,0,0) fanout_n_80 (N373, {N373_0, N373_1});
fanout_n #(2,0,0) fanout_n_81 (N376, {N376_0, N376_1});
fanout_n #(2,0,0) fanout_n_82 (N379, {N379_0, N379_1});
fanout_n #(2,0,0) fanout_n_83 (N382, {N382_0, N382_1});
fanout_n #(2,0,0) fanout_n_84 (N385, {N385_0, N385_1});
fanout_n #(2,0,0) fanout_n_85 (N388, {N388_0, N388_1});
fanout_n #(2,0,0) fanout_n_86 (N556, {N556_0, N556_1});
fanout_n #(2,0,0) fanout_n_87 (N559, {N559_0, N559_1});
fanout_n #(2,0,0) fanout_n_88 (N562, {N562_0, N562_1});
fanout_n #(2,0,0) fanout_n_89 (N565, {N565_0, N565_1});
fanout_n #(2,0,0) fanout_n_90 (N568, {N568_0, N568_1});
fanout_n #(2,0,0) fanout_n_91 (N571, {N571_0, N571_1});
fanout_n #(2,0,0) fanout_n_92 (N574, {N574_0, N574_1});
fanout_n #(2,0,0) fanout_n_93 (N577, {N577_0, N577_1});
fanout_n #(2,0,0) fanout_n_94 (N580, {N580_0, N580_1});
fanout_n #(2,0,0) fanout_n_95 (N583, {N583_0, N583_1});
fanout_n #(2,0,0) fanout_n_96 (N586, {N586_0, N586_1});
fanout_n #(2,0,0) fanout_n_97 (N589, {N589_0, N589_1});
fanout_n #(2,0,0) fanout_n_98 (N592, {N592_0, N592_1});
fanout_n #(2,0,0) fanout_n_99 (N595, {N595_0, N595_1});
fanout_n #(2,0,0) fanout_n_100 (N598, {N598_0, N598_1});
fanout_n #(4,0,0) fanout_n_101 (N603, {N603_0, N603_1, N603_2, N603_3});
fanout_n #(3,0,0) fanout_n_102 (N608, {N608_0, N608_1, N608_2});
fanout_n #(3,0,0) fanout_n_103 (N612, {N612_0, N612_1, N612_2});
fanout_n #(2,0,0) fanout_n_104 (N616, {N616_0, N616_1});
fanout_n #(2,0,0) fanout_n_105 (N619, {N619_0, N619_1});
fanout_n #(2,0,0) fanout_n_106 (N622, {N622_0, N622_1});
fanout_n #(2,0,0) fanout_n_107 (N625, {N625_0, N625_1});
fanout_n #(2,0,0) fanout_n_108 (N628, {N628_0, N628_1});
fanout_n #(2,0,0) fanout_n_109 (N631, {N631_0, N631_1});
fanout_n #(2,0,0) fanout_n_110 (N634, {N634_0, N634_1});
fanout_n #(2,0,0) fanout_n_111 (N637, {N637_0, N637_1});
fanout_n #(2,0,0) fanout_n_112 (N640, {N640_0, N640_1});
fanout_n #(2,0,0) fanout_n_113 (N643, {N643_0, N643_1});
fanout_n #(2,0,0) fanout_n_114 (N646, {N646_0, N646_1});
fanout_n #(2,0,0) fanout_n_115 (N649, {N649_0, N649_1});
fanout_n #(2,0,0) fanout_n_116 (N652, {N652_0, N652_1});
fanout_n #(2,0,0) fanout_n_117 (N655, {N655_0, N655_1});
fanout_n #(2,0,0) fanout_n_118 (N658, {N658_0, N658_1});
fanout_n #(2,0,0) fanout_n_119 (N661, {N661_0, N661_1});
fanout_n #(2,0,0) fanout_n_120 (N664, {N664_0, N664_1});
fanout_n #(2,0,0) fanout_n_121 (N667, {N667_0, N667_1});
fanout_n #(2,0,0) fanout_n_122 (N670, {N670_0, N670_1});
fanout_n #(2,0,0) fanout_n_123 (N673, {N673_0, N673_1});
fanout_n #(2,0,0) fanout_n_124 (N676, {N676_0, N676_1});
fanout_n #(2,0,0) fanout_n_125 (N679, {N679_0, N679_1});
fanout_n #(2,0,0) fanout_n_126 (N682, {N682_0, N682_1});
fanout_n #(2,0,0) fanout_n_127 (N685, {N685_0, N685_1});
fanout_n #(2,0,0) fanout_n_128 (N688, {N688_0, N688_1});
fanout_n #(2,0,0) fanout_n_129 (N691, {N691_0, N691_1});
fanout_n #(2,0,0) fanout_n_130 (N694, {N694_0, N694_1});
fanout_n #(2,0,0) fanout_n_131 (N697, {N697_0, N697_1});
fanout_n #(2,0,0) fanout_n_132 (N700, {N700_0, N700_1});
fanout_n #(2,0,0) fanout_n_133 (N703, {N703_0, N703_1});
fanout_n #(2,0,0) fanout_n_134 (N706, {N706_0, N706_1});
fanout_n #(2,0,0) fanout_n_135 (N709, {N709_0, N709_1});
fanout_n #(2,0,0) fanout_n_136 (N712, {N712_0, N712_1});
fanout_n #(2,0,0) fanout_n_137 (N715, {N715_0, N715_1});
fanout_n #(2,0,0) fanout_n_138 (N718, {N718_0, N718_1});
fanout_n #(2,0,0) fanout_n_139 (N721, {N721_0, N721_1});
fanout_n #(2,0,0) fanout_n_140 (N724, {N724_0, N724_1});
fanout_n #(2,0,0) fanout_n_141 (N727, {N727_0, N727_1});
fanout_n #(2,0,0) fanout_n_142 (N730, {N730_0, N730_1});
fanout_n #(2,0,0) fanout_n_143 (N733, {N733_0, N733_1});
fanout_n #(2,0,0) fanout_n_144 (N736, {N736_0, N736_1});
fanout_n #(2,0,0) fanout_n_145 (N739, {N739_0, N739_1});
fanout_n #(2,0,0) fanout_n_146 (N742, {N742_0, N742_1});
fanout_n #(2,0,0) fanout_n_147 (N745, {N745_0, N745_1});
fanout_n #(2,0,0) fanout_n_148 (N748, {N748_0, N748_1});
fanout_n #(2,0,0) fanout_n_149 (N751, {N751_0, N751_1});
fanout_n #(3,0,0) fanout_n_150 (N899, {N899_0, N899_1, N899_2});
fanout_n #(3,0,0) fanout_n_151 (N903, {N903_0, N903_1, N903_2});
fanout_n #(2,0,0) fanout_n_152 (N907, {N907_0, N907_1});
fanout_n #(2,0,0) fanout_n_153 (N910, {N910_0, N910_1});
fanout_n #(2,0,0) fanout_n_154 (N923, {N923_0, N923_1});
fanout_n #(8,0,0) fanout_n_155 (N926, {N926_0, N926_1, N926_2, N926_3, N926_4, N926_5, N926_6, N926_7});
fanout_n #(2,0,0) fanout_n_156 (N935, {N935_0, N935_1});
fanout_n #(2,0,0) fanout_n_157 (N939, {N939_0, N939_1});
fanout_n #(2,0,0) fanout_n_158 (N943, {N943_0, N943_1});
fanout_n #(2,0,0) fanout_n_159 (N947, {N947_0, N947_1});
fanout_n #(2,0,0) fanout_n_160 (N951, {N951_0, N951_1});
fanout_n #(2,0,0) fanout_n_161 (N955, {N955_0, N955_1});
fanout_n #(2,0,0) fanout_n_162 (N959, {N959_0, N959_1});
fanout_n #(2,0,0) fanout_n_163 (N962, {N962_0, N962_1});
fanout_n #(2,0,0) fanout_n_164 (N965, {N965_0, N965_1});
fanout_n #(2,0,0) fanout_n_165 (N969, {N969_0, N969_1});
fanout_n #(2,0,0) fanout_n_166 (N973, {N973_0, N973_1});
fanout_n #(2,0,0) fanout_n_167 (N977, {N977_0, N977_1});
fanout_n #(2,0,0) fanout_n_168 (N981, {N981_0, N981_1});
fanout_n #(2,0,0) fanout_n_169 (N985, {N985_0, N985_1});
fanout_n #(2,0,0) fanout_n_170 (N994, {N994_0, N994_1});
fanout_n #(2,0,0) fanout_n_171 (N998, {N998_0, N998_1});
fanout_n #(2,0,0) fanout_n_172 (N1010, {N1010_0, N1010_1});
fanout_n #(2,0,0) fanout_n_173 (N1013, {N1013_0, N1013_1});
fanout_n #(2,0,0) fanout_n_174 (N1016, {N1016_0, N1016_1});
fanout_n #(2,0,0) fanout_n_175 (N1019, {N1019_0, N1019_1});
fanout_n #(2,0,0) fanout_n_176 (N1022, {N1022_0, N1022_1});
fanout_n #(2,0,0) fanout_n_177 (N1025, {N1025_0, N1025_1});
fanout_n #(2,0,0) fanout_n_178 (N1028, {N1028_0, N1028_1});
fanout_n #(2,0,0) fanout_n_179 (N1031, {N1031_0, N1031_1});
fanout_n #(2,0,0) fanout_n_180 (N1034, {N1034_0, N1034_1});
fanout_n #(2,0,0) fanout_n_181 (N1037, {N1037_0, N1037_1});
fanout_n #(2,0,0) fanout_n_182 (N1040, {N1040_0, N1040_1});
fanout_n #(2,0,0) fanout_n_183 (N1043, {N1043_0, N1043_1});
fanout_n #(2,0,0) fanout_n_184 (N1046, {N1046_0, N1046_1});
fanout_n #(2,0,0) fanout_n_185 (N1049, {N1049_0, N1049_1});
fanout_n #(2,0,0) fanout_n_186 (N1164, {N1164_0, N1164_1});
fanout_n #(2,0,0) fanout_n_187 (N1168, {N1168_0, N1168_1});
fanout_n #(16,0,0) fanout_n_188 (N1171, {N1171_0, N1171_1, N1171_2, N1171_3, N1171_4, N1171_5, N1171_6, N1171_7, N1171_8, N1171_9, N1171_10, N1171_11, N1171_12, N1171_13, N1171_14, N1171_15});
fanout_n #(16,0,0) fanout_n_189 (N1188, {N1188_0, N1188_1, N1188_2, N1188_3, N1188_4, N1188_5, N1188_6, N1188_7, N1188_8, N1188_9, N1188_10, N1188_11, N1188_12, N1188_13, N1188_14, N1188_15});
fanout_n #(2,0,0) fanout_n_190 (N1232, {N1232_0, N1232_1});
fanout_n #(2,0,0) fanout_n_191 (N1235, {N1235_0, N1235_1});
fanout_n #(2,0,0) fanout_n_192 (N1243, {N1243_0, N1243_1});
fanout_n #(2,0,0) fanout_n_193 (N1246, {N1246_0, N1246_1});
fanout_n #(2,0,0) fanout_n_194 (N1249, {N1249_0, N1249_1});
fanout_n #(2,0,0) fanout_n_195 (N1252, {N1252_0, N1252_1});
fanout_n #(2,0,0) fanout_n_196 (N1255, {N1255_0, N1255_1});
fanout_n #(2,0,0) fanout_n_197 (N1258, {N1258_0, N1258_1});
fanout_n #(2,0,0) fanout_n_198 (N1261, {N1261_0, N1261_1});
fanout_n #(2,0,0) fanout_n_199 (N1264, {N1264_0, N1264_1});
fanout_n #(2,0,0) fanout_n_200 (N1319, {N1319_0, N1319_1});
fanout_n #(2,0,0) fanout_n_201 (N1334, {N1334_0, N1334_1});
fanout_n #(2,0,0) fanout_n_202 (N1352, {N1352_0, N1352_1});
fanout_n #(2,0,0) fanout_n_203 (N1355, {N1355_0, N1355_1});
fanout_n #(2,0,0) fanout_n_204 (N1358, {N1358_0, N1358_1});
fanout_n #(2,0,0) fanout_n_205 (N1361, {N1361_0, N1361_1});
fanout_n #(2,0,0) fanout_n_206 (N1364, {N1364_0, N1364_1});
fanout_n #(2,0,0) fanout_n_207 (N1367, {N1367_0, N1367_1});
fanout_n #(2,0,0) fanout_n_208 (N1370, {N1370_0, N1370_1});
fanout_n #(2,0,0) fanout_n_209 (N1373, {N1373_0, N1373_1});
fanout_n #(2,0,0) fanout_n_210 (N1376, {N1376_0, N1376_1});
fanout_n #(2,0,0) fanout_n_211 (N1379, {N1379_0, N1379_1});
fanout_n #(2,0,0) fanout_n_212 (N1383, {N1383_0, N1383_1});
fanout_n #(2,0,0) fanout_n_213 (N1390, {N1390_0, N1390_1});
fanout_n #(2,0,0) fanout_n_214 (N1393, {N1393_0, N1393_1});
fanout_n #(2,0,0) fanout_n_215 (N1416, {N1416_0, N1416_1});
fanout_n #(2,0,0) fanout_n_216 (N1419, {N1419_0, N1419_1});
fanout_n #(2,0,0) fanout_n_217 (N1440, {N1440_0, N1440_1});
fanout_n #(2,0,0) fanout_n_218 (N1472, {N1472_0, N1472_1});
fanout_n #(2,0,0) fanout_n_219 (N1478, {N1478_0, N1478_1});
fanout_n #(2,0,0) fanout_n_220 (N1481, {N1481_0, N1481_1});
fanout_n #(2,0,0) fanout_n_221 (N1484, {N1484_0, N1484_1});
fanout_n #(2,0,0) fanout_n_222 (N1510, {N1510_0, N1510_1});
fanout_n #(2,0,0) fanout_n_223 (N1514, {N1514_0, N1514_1});
fanout_n #(2,0,0) fanout_n_224 (N1517, {N1517_0, N1517_1});
fanout_n #(3,0,0) fanout_n_225 (N1522, {N1522_0, N1522_1, N1522_2});
fanout_n #(2,0,0) fanout_n_226 (N1534, {N1534_0, N1534_1});
fanout_n #(2,0,0) fanout_n_227 (N1537, {N1537_0, N1537_1});
fanout_n #(2,0,0) fanout_n_228 (N1540, {N1540_0, N1540_1});
fanout_n #(2,0,0) fanout_n_229 (N1546, {N1546_0, N1546_1});
fanout_n #(2,0,0) fanout_n_230 (N1554, {N1554_0, N1554_1});
fanout_n #(3,0,0) fanout_n_231 (N1557, {N1557_0, N1557_1, N1557_2});
fanout_n #(2,0,0) fanout_n_232 (N1561, {N1561_0, N1561_1});
fanout_n #(2,0,0) fanout_n_233 (N1571, {N1571_0, N1571_1});
fanout_n #(2,0,0) fanout_n_234 (N1576, {N1576_0, N1576_1});
fanout_n #(2,0,0) fanout_n_235 (N1588, {N1588_0, N1588_1});
fanout_n #(2,0,0) fanout_n_236 (N1596, {N1596_0, N1596_1});
fanout_n #(2,0,0) fanout_n_237 (N1600, {N1600_0, N1600_1});
fanout_n #(2,0,0) fanout_n_238 (N1603, {N1603_0, N1603_1});
fanout_n #(2,0,0) fanout_n_239 (N1606, {N1606_0, N1606_1});
fanout_n #(2,0,0) fanout_n_240 (N1609, {N1609_0, N1609_1});
fanout_n #(2,0,0) fanout_n_241 (N1612, {N1612_0, N1612_1});
fanout_n #(2,0,0) fanout_n_242 (N1615, {N1615_0, N1615_1});
fanout_n #(2,0,0) fanout_n_243 (N1620, {N1620_0, N1620_1});
fanout_n #(2,0,0) fanout_n_244 (N1623, {N1623_0, N1623_1});
fanout_n #(2,0,0) fanout_n_245 (N1640, {N1640_0, N1640_1});
fanout_n #(2,0,0) fanout_n_246 (N1643, {N1643_0, N1643_1});
fanout_n #(2,0,0) fanout_n_247 (N1647, {N1647_0, N1647_1});
fanout_n #(2,0,0) fanout_n_248 (N1651, {N1651_0, N1651_1});
fanout_n #(2,0,0) fanout_n_249 (N1658, {N1658_0, N1658_1});
fanout_n #(2,0,0) fanout_n_250 (N1661, {N1661_0, N1661_1});
fanout_n #(2,0,0) fanout_n_251 (N1664, {N1664_0, N1664_1});
fanout_n #(2,0,0) fanout_n_252 (N1685, {N1685_0, N1685_1});
fanout_n #(2,0,0) fanout_n_253 (N1697, {N1697_0, N1697_1});
fanout_n #(2,0,0) fanout_n_254 (N1701, {N1701_0, N1701_1});
fanout_n #(2,0,0) fanout_n_255 (N1714, {N1714_0, N1714_1});
fanout_n #(2,0,0) fanout_n_256 (N1717, {N1717_0, N1717_1});
fanout_n #(2,0,0) fanout_n_257 (N1723, {N1723_0, N1723_1});
fanout_n #(2,0,0) fanout_n_258 (N1731, {N1731_0, N1731_1});
fanout_n #(2,0,0) fanout_n_259 (N1734, {N1734_0, N1734_1});
fanout_n #(2,0,0) fanout_n_260 (N1742, {N1742_0, N1742_1});
fanout_n #(2,0,0) fanout_n_261 (N1748, {N1748_0, N1748_1});
fanout_n #(2,0,0) fanout_n_262 (N1751, {N1751_0, N1751_1});
fanout_n #(2,0,0) fanout_n_263 (N1774, {N1774_0, N1774_1});
fanout_n #(2,0,0) fanout_n_264 (N1777, {N1777_0, N1777_1});
fanout_n #(2,0,0) fanout_n_265 (N1788, {N1788_0, N1788_1});
fanout_n #(2,0,0) fanout_n_266 (N1798, {N1798_0, N1798_1});
fanout_n #(2,0,0) fanout_n_267 (N1802, {N1802_0, N1802_1});
fanout_n #(2,0,0) fanout_n_268 (N1812, {N1812_0, N1812_1});
fanout_n #(2,0,0) fanout_n_269 (N1815, {N1815_0, N1815_1});
fanout_n #(2,0,0) fanout_n_270 (N1818, {N1818_0, N1818_1});
fanout_n #(2,0,0) fanout_n_271 (N1830, {N1830_0, N1830_1});
fanout_n #(2,0,0) fanout_n_272 (N1838, {N1838_0, N1838_1});
fanout_n #(2,0,0) fanout_n_273 (N1841, {N1841_0, N1841_1});
fanout_n #(2,0,0) fanout_n_274 (N1858, {N1858_0, N1858_1});
fanout_n #(2,0,0) fanout_n_275 (N1866, {N1866_0, N1866_1});
fanout_n #(2,0,0) fanout_n_276 (N1869, {N1869_0, N1869_1});
fanout_n #(2,0,0) fanout_n_277 (N1872, {N1872_0, N1872_1});
fanout_n #(2,0,0) fanout_n_278 (N1875, {N1875_0, N1875_1});
fanout_n #(2,0,0) fanout_n_279 (N1879, {N1879_0, N1879_1});
fanout_n #(2,0,0) fanout_n_280 (N1889, {N1889_0, N1889_1});
fanout_n #(2,0,0) fanout_n_281 (N1898, {N1898_0, N1898_1});
fanout_n #(2,0,0) fanout_n_282 (N1902, {N1902_0, N1902_1});
fanout_n #(2,0,0) fanout_n_283 (N1927, {N1927_0, N1927_1});
fanout_n #(2,0,0) fanout_n_284 (N1930, {N1930_0, N1930_1});
fanout_n #(2,0,0) fanout_n_285 (N1933, {N1933_0, N1933_1});
fanout_n #(2,0,0) fanout_n_286 (N1944, {N1944_0, N1944_1});
fanout_n #(2,0,0) fanout_n_287 (N1947, {N1947_0, N1947_1});
fanout_n #(2,0,0) fanout_n_288 (N1950, {N1950_0, N1950_1});
fanout_n #(2,0,0) fanout_n_289 (N1953, {N1953_0, N1953_1});
fanout_n #(2,0,0) fanout_n_290 (N1958, {N1958_0, N1958_1});
fanout_n #(2,0,0) fanout_n_291 (N1961, {N1961_0, N1961_1});
fanout_n #(2,0,0) fanout_n_292 (N1965, {N1965_0, N1965_1});
fanout_n #(2,0,0) fanout_n_293 (N1968, {N1968_0, N1968_1});
fanout_n #(2,0,0) fanout_n_294 (N1980, {N1980_0, N1980_1});
fanout_n #(2,0,0) fanout_n_295 (N1987, {N1987_0, N1987_1});
fanout_n #(2,0,0) fanout_n_296 (N2027, {N2027_0, N2027_1});
fanout_n #(2,0,0) fanout_n_297 (N2030, {N2030_0, N2030_1});
fanout_n #(2,0,0) fanout_n_298 (N2033, {N2033_0, N2033_1});
fanout_n #(2,0,0) fanout_n_299 (N2042, {N2042_0, N2042_1});
fanout_n #(2,0,0) fanout_n_300 (N2052, {N2052_0, N2052_1});
fanout_n #(2,0,0) fanout_n_301 (N2055, {N2055_0, N2055_1});
fanout_n #(2,0,0) fanout_n_302 (N2062, {N2062_0, N2062_1});
fanout_n #(2,0,0) fanout_n_303 (N2068, {N2068_0, N2068_1});
fanout_n #(2,0,0) fanout_n_304 (N2071, {N2071_0, N2071_1});
fanout_n #(2,0,0) fanout_n_305 (N2078, {N2078_0, N2078_1});
fanout_n #(2,0,0) fanout_n_306 (N2081, {N2081_0, N2081_1});
fanout_n #(2,0,0) fanout_n_307 (N2086, {N2086_0, N2086_1});
fanout_n #(2,0,0) fanout_n_308 (N2089, {N2089_0, N2089_1});
fanout_n #(14,0,0) fanout_n_309 (N2104, {N2104_0, N2104_1, N2104_2, N2104_3, N2104_4, N2104_5, N2104_6, N2104_7, N2104_8, N2104_9, N2104_10, N2104_11, N2104_12, N2104_13});
fanout_n #(9,0,0) fanout_n_310 (N2119, {N2119_0, N2119_1, N2119_2, N2119_3, N2119_4, N2119_5, N2119_6, N2119_7, N2119_8});
fanout_n #(13,0,0) fanout_n_311 (N2129, {N2129_0, N2129_1, N2129_2, N2129_3, N2129_4, N2129_5, N2129_6, N2129_7, N2129_8, N2129_9, N2129_10, N2129_11, N2129_12});
fanout_n #(4,0,0) fanout_n_312 (N2143, {N2143_0, N2143_1, N2143_2, N2143_3});
fanout_n #(2,0,0) fanout_n_313 (N2148, {N2148_0, N2148_1});
fanout_n #(2,0,0) fanout_n_314 (N2151, {N2151_0, N2151_1});
fanout_n #(2,0,0) fanout_n_315 (N2196, {N2196_0, N2196_1});
fanout_n #(2,0,0) fanout_n_316 (N2199, {N2199_0, N2199_1});
fanout_n #(2,0,0) fanout_n_317 (N2202, {N2202_0, N2202_1});
fanout_n #(2,0,0) fanout_n_318 (N2205, {N2205_0, N2205_1});
fanout_n #(2,0,0) fanout_n_319 (N2237, {N2237_0, N2237_1});
fanout_n #(2,0,0) fanout_n_320 (N2241, {N2241_0, N2241_1});
fanout_n #(2,0,0) fanout_n_321 (N2245, {N2245_0, N2245_1});
fanout_n #(2,0,0) fanout_n_322 (N2257, {N2257_0, N2257_1});
fanout_n #(2,0,0) fanout_n_323 (N2260, {N2260_0, N2260_1});
fanout_n #(2,0,0) fanout_n_324 (N2263, {N2263_0, N2263_1});
fanout_n #(2,0,0) fanout_n_325 (N2266, {N2266_0, N2266_1});
fanout_n #(2,0,0) fanout_n_326 (N2269, {N2269_0, N2269_1});
fanout_n #(2,0,0) fanout_n_327 (N2272, {N2272_0, N2272_1});
fanout_n #(2,0,0) fanout_n_328 (N2279, {N2279_0, N2279_1});
fanout_n #(10,0,0) fanout_n_329 (N2286, {N2286_0, N2286_1, N2286_2, N2286_3, N2286_4, N2286_5, N2286_6, N2286_7, N2286_8, N2286_9});
fanout_n #(15,0,0) fanout_n_330 (N2297, {N2297_0, N2297_1, N2297_2, N2297_3, N2297_4, N2297_5, N2297_6, N2297_7, N2297_8, N2297_9, N2297_10, N2297_11, N2297_12, N2297_13, N2297_14});
fanout_n #(10,0,0) fanout_n_331 (N2315, {N2315_0, N2315_1, N2315_2, N2315_3, N2315_4, N2315_5, N2315_6, N2315_7, N2315_8, N2315_9});
fanout_n #(13,0,0) fanout_n_332 (N2326, {N2326_0, N2326_1, N2326_2, N2326_3, N2326_4, N2326_5, N2326_6, N2326_7, N2326_8, N2326_9, N2326_10, N2326_11, N2326_12});
fanout_n #(12,0,0) fanout_n_333 (N2340, {N2340_0, N2340_1, N2340_2, N2340_3, N2340_4, N2340_5, N2340_6, N2340_7, N2340_8, N2340_9, N2340_10, N2340_11});
fanout_n #(7,0,0) fanout_n_334 (N2353, {N2353_0, N2353_1, N2353_2, N2353_3, N2353_4, N2353_5, N2353_6});
fanout_n #(13,0,0) fanout_n_335 (N2361, {N2361_0, N2361_1, N2361_2, N2361_3, N2361_4, N2361_5, N2361_6, N2361_7, N2361_8, N2361_9, N2361_10, N2361_11, N2361_12});
fanout_n #(8,0,0) fanout_n_336 (N2375, {N2375_0, N2375_1, N2375_2, N2375_3, N2375_4, N2375_5, N2375_6, N2375_7});
fanout_n #(14,0,0) fanout_n_337 (N2386, {N2386_0, N2386_1, N2386_2, N2386_3, N2386_4, N2386_5, N2386_6, N2386_7, N2386_8, N2386_9, N2386_10, N2386_11, N2386_12, N2386_13});
fanout_n #(16,0,0) fanout_n_338 (N2427, {N2427_0, N2427_1, N2427_2, N2427_3, N2427_4, N2427_5, N2427_6, N2427_7, N2427_8, N2427_9, N2427_10, N2427_11, N2427_12, N2427_13, N2427_14, N2427_15});
fanout_n #(2,0,0) fanout_n_339 (N2537, {N2537_0, N2537_1});
fanout_n #(2,0,0) fanout_n_340 (N2540, {N2540_0, N2540_1});
fanout_n #(2,0,0) fanout_n_341 (N2543, {N2543_0, N2543_1});
fanout_n #(2,0,0) fanout_n_342 (N2546, {N2546_0, N2546_1});
fanout_n #(2,0,0) fanout_n_343 (N2549, {N2549_0, N2549_1});
fanout_n #(2,0,0) fanout_n_344 (N2552, {N2552_0, N2552_1});
fanout_n #(2,0,0) fanout_n_345 (N2555, {N2555_0, N2555_1});
fanout_n #(2,0,0) fanout_n_346 (N2558, {N2558_0, N2558_1});
fanout_n #(2,0,0) fanout_n_347 (N2561, {N2561_0, N2561_1});
fanout_n #(2,0,0) fanout_n_348 (N2564, {N2564_0, N2564_1});
fanout_n #(2,0,0) fanout_n_349 (N2567, {N2567_0, N2567_1});
fanout_n #(2,0,0) fanout_n_350 (N2570, {N2570_0, N2570_1});
fanout_n #(2,0,0) fanout_n_351 (N2573, {N2573_0, N2573_1});
fanout_n #(2,0,0) fanout_n_352 (N2576, {N2576_0, N2576_1});
fanout_n #(2,0,0) fanout_n_353 (N2594, {N2594_0, N2594_1});
fanout_n #(2,0,0) fanout_n_354 (N2597, {N2597_0, N2597_1});
fanout_n #(2,0,0) fanout_n_355 (N2600, {N2600_0, N2600_1});
fanout_n #(2,0,0) fanout_n_356 (N2603, {N2603_0, N2603_1});
fanout_n #(2,0,0) fanout_n_357 (N2606, {N2606_0, N2606_1});
fanout_n #(2,0,0) fanout_n_358 (N2611, {N2611_0, N2611_1});
fanout_n #(2,0,0) fanout_n_359 (N2614, {N2614_0, N2614_1});
fanout_n #(2,0,0) fanout_n_360 (N2617, {N2617_0, N2617_1});
fanout_n #(2,0,0) fanout_n_361 (N2620, {N2620_0, N2620_1});
fanout_n #(2,0,0) fanout_n_362 (N2639, {N2639_0, N2639_1});
fanout_n #(2,0,0) fanout_n_363 (N2642, {N2642_0, N2642_1});
fanout_n #(2,0,0) fanout_n_364 (N2645, {N2645_0, N2645_1});
fanout_n #(2,0,0) fanout_n_365 (N2648, {N2648_0, N2648_1});
fanout_n #(2,0,0) fanout_n_366 (N2651, {N2651_0, N2651_1});
fanout_n #(2,0,0) fanout_n_367 (N2655, {N2655_0, N2655_1});
fanout_n #(2,0,0) fanout_n_368 (N2658, {N2658_0, N2658_1});
fanout_n #(2,0,0) fanout_n_369 (N2661, {N2661_0, N2661_1});
fanout_n #(2,0,0) fanout_n_370 (N2664, {N2664_0, N2664_1});
fanout_n #(2,0,0) fanout_n_371 (N2747, {N2747_0, N2747_1});
fanout_n #(2,0,0) fanout_n_372 (N2750, {N2750_0, N2750_1});
fanout_n #(2,0,0) fanout_n_373 (N2773, {N2773_0, N2773_1});
fanout_n #(2,0,0) fanout_n_374 (N2776, {N2776_0, N2776_1});
fanout_n #(6,0,0) fanout_n_375 (N2789, {N2789_0, N2789_1, N2789_2, N2789_3, N2789_4, N2789_5});
fanout_n #(2,0,0) fanout_n_376 (N2812, {N2812_0, N2812_1});
fanout_n #(2,0,0) fanout_n_377 (N2815, {N2815_0, N2815_1});
fanout_n #(2,0,0) fanout_n_378 (N2818, {N2818_0, N2818_1});
fanout_n #(2,0,0) fanout_n_379 (N2821, {N2821_0, N2821_1});
fanout_n #(2,0,0) fanout_n_380 (N2824, {N2824_0, N2824_1});
fanout_n #(2,0,0) fanout_n_381 (N2829, {N2829_0, N2829_1});
fanout_n #(2,0,0) fanout_n_382 (N2843, {N2843_0, N2843_1});
fanout_n #(2,0,0) fanout_n_383 (N2846, {N2846_0, N2846_1});
fanout_n #(2,0,0) fanout_n_384 (N2883, {N2883_0, N2883_1});


notg NOT1_1 (N190, N1_0);
notg NOT1_2 (N194, N4_0);
notg NOT1_3 (N197, N7_0);
notg NOT1_4 (N201, N10_0);
notg NOT1_5 (N206, N13_0);
notg NOT1_6 (N209, N16_0);
notg NOT1_7 (N212, N19_0);
notg NOT1_8 (N216, N22_0);
notg NOT1_9 (N220, N25_0);
notg NOT1_10 (N225, N28_0);
notg NOT1_11 (N229, N31_0);
notg NOT1_12 (N232, N34_0);
notg NOT1_13 (N235, N37_0);
notg NOT1_14 (N239, N40_0);
notg NOT1_15 (N243, N43_0);
notg NOT1_16 (N247, N46_0);
nand_n #(2,0,0) NAND2_17 (N251, {N63_0, N88_0});
nand_n #(2,0,0) NAND2_18 (N252, {N66_0, N91_0});
notg NOT1_19 (N253, N72_0);
notg NOT1_20 (N256, N72_1);
bufg BUFF1_21 (N257, N69_0);
bufg BUFF1_22 (N260, N69_1);
notg NOT1_23 (N263, N76_0);
notg NOT1_24 (N266, N79_0);
notg NOT1_25 (N269, N82_0);
notg NOT1_26 (N272, N85_0);
notg NOT1_27 (N275, N104_0);
notg NOT1_28 (N276, N104_1);
notg NOT1_29 (N277, N88_1);
notg NOT1_30 (N280, N91_1);
bufg BUFF1_31 (N283, N94_0);
notg NOT1_32 (N290, N94_1);
bufg BUFF1_33 (N297, N94_2);
notg NOT1_34 (N300, N94_3);
bufg BUFF1_35 (N303, N99_0);
notg NOT1_36 (N306, N99_1);
notg NOT1_37 (N313, N99_2);
bufg BUFF1_38 (N316, N104_2);
notg NOT1_39 (N319, N104_3);
bufg BUFF1_40 (N326, N104_4);
bufg BUFF1_41 (N331, N104_5);
notg NOT1_42 (N338, N104_6);
bufg BUFF1_43 (N343, N1_1);
bufg BUFF1_44 (N346, N4_1);
bufg BUFF1_45 (N349, N7_1);
bufg BUFF1_46 (N352, N10_1);
bufg BUFF1_47 (N355, N13_1);
bufg BUFF1_48 (N358, N16_1);
bufg BUFF1_49 (N361, N19_1);
bufg BUFF1_50 (N364, N22_1);
bufg BUFF1_51 (N367, N25_1);
bufg BUFF1_52 (N370, N28_1);
bufg BUFF1_53 (N373, N31_1);
bufg BUFF1_54 (N376, N34_1);
bufg BUFF1_55 (N379, N37_1);
bufg BUFF1_56 (N382, N40_1);
bufg BUFF1_57 (N385, N43_1);
bufg BUFF1_58 (N388, N46_1);
notg NOT1_59 (N534, N343_0);
notg NOT1_60 (N535, N346_0);
notg NOT1_61 (N536, N349_0);
notg NOT1_62 (N537, N352_0);
notg NOT1_63 (N538, N355_0);
notg NOT1_64 (N539, N358_0);
notg NOT1_65 (N540, N361_0);
notg NOT1_66 (N541, N364_0);
notg NOT1_67 (N542, N367_0);
notg NOT1_68 (N543, N370_0);
notg NOT1_69 (N544, N373_0);
notg NOT1_70 (N545, N376_0);
notg NOT1_71 (N546, N379_0);
notg NOT1_72 (N547, N382_0);
notg NOT1_73 (N548, N385_0);
notg NOT1_74 (N549, N388_0);
nand_n #(2,0,0) NAND2_75 (N550, {N306_0, N331_0});
nand_n #(2,0,0) NAND2_76 (N551, {N306_1, N331_1});
nand_n #(2,0,0) NAND2_77 (N552, {N306_2, N331_2});
nand_n #(2,0,0) NAND2_78 (N553, {N306_3, N331_3});
nand_n #(2,0,0) NAND2_79 (N554, {N306_4, N331_4});
nand_n #(2,0,0) NAND2_80 (N555, {N306_5, N331_5});
bufg BUFF1_81 (N556, N190_0);
bufg BUFF1_82 (N559, N194_0);
bufg BUFF1_83 (N562, N206_0);
bufg BUFF1_84 (N565, N209_0);
bufg BUFF1_85 (N568, N225_0);
bufg BUFF1_86 (N571, N243_0);
and_n #(2,0,0) AND2_87 (N574, {N63_1, N319_0});
bufg BUFF1_88 (N577, N220_0);
bufg BUFF1_89 (N580, N229_0);
bufg BUFF1_90 (N583, N232_0);
and_n #(2,0,0) AND2_91 (N586, {N66_1, N319_1});
bufg BUFF1_92 (N589, N239_0);
and_n #(3,0,0) AND3_93 (N592, {N49_0, N253_0, N319_2});
bufg BUFF1_94 (N595, N247_0);
bufg BUFF1_95 (N598, N239_1);
nand_n #(2,0,0) NAND2_96 (N601, {N326_0, N277_0});
nand_n #(2,0,0) NAND2_97 (N602, {N326_1, N280_0});
nand_n #(2,0,0) NAND2_98 (N603, {N260_0, N72_2});
nand_n #(2,0,0) NAND2_99 (N608, {N260_1, N300_0});
nand_n #(2,0,0) NAND2_100 (N612, {N256, N300_1});
bufg BUFF1_101 (N616, N201_0);
bufg BUFF1_102 (N619, N216_0);
bufg BUFF1_103 (N622, N220_1);
bufg BUFF1_104 (N625, N239_2);
bufg BUFF1_105 (N628, N190_1);
bufg BUFF1_106 (N631, N190_2);
bufg BUFF1_107 (N634, N194_1);
bufg BUFF1_108 (N637, N229_1);
bufg BUFF1_109 (N640, N197_0);
and_n #(3,0,0) AND3_110 (N643, {N56_0, N257_0, N319_3});
bufg BUFF1_111 (N646, N232_1);
bufg BUFF1_112 (N649, N201_1);
bufg BUFF1_113 (N652, N235_0);
and_n #(3,0,0) AND3_114 (N655, {N60_0, N257_1, N319_4});
bufg BUFF1_115 (N658, N263_0);
bufg BUFF1_116 (N661, N263_1);
bufg BUFF1_117 (N664, N266_0);
bufg BUFF1_118 (N667, N266_1);
bufg BUFF1_119 (N670, N269_0);
bufg BUFF1_120 (N673, N269_1);
bufg BUFF1_121 (N676, N272_0);
bufg BUFF1_122 (N679, N272_1);
and_n #(2,0,0) AND2_123 (N682, {N251, N316_0});
and_n #(2,0,0) AND2_124 (N685, {N252, N316_1});
bufg BUFF1_125 (N688, N197_1);
bufg BUFF1_126 (N691, N197_2);
bufg BUFF1_127 (N694, N212_0);
bufg BUFF1_128 (N697, N212_1);
bufg BUFF1_129 (N700, N247_1);
bufg BUFF1_130 (N703, N247_2);
bufg BUFF1_131 (N706, N235_1);
bufg BUFF1_132 (N709, N235_2);
bufg BUFF1_133 (N712, N201_2);
bufg BUFF1_134 (N715, N201_3);
bufg BUFF1_135 (N718, N206_1);
bufg BUFF1_136 (N721, N216_1);
and_n #(3,0,0) AND3_137 (N724, {N53_0, N253_1, N319_5});
bufg BUFF1_138 (N727, N243_1);
bufg BUFF1_139 (N730, N220_2);
bufg BUFF1_140 (N733, N220_3);
bufg BUFF1_141 (N736, N209_1);
bufg BUFF1_142 (N739, N216_2);
bufg BUFF1_143 (N742, N225_1);
bufg BUFF1_144 (N745, N243_2);
bufg BUFF1_145 (N748, N212_2);
bufg BUFF1_146 (N751, N225_2);
notg NOT1_147 (N886, N682_0);
notg NOT1_148 (N887, N685_0);
notg NOT1_149 (N888, N616_0);
notg NOT1_150 (N889, N619_0);
notg NOT1_151 (N890, N622_0);
notg NOT1_152 (N891, N625_0);
notg NOT1_153 (N892, N631_0);
notg NOT1_154 (N893, N643_0);
notg NOT1_155 (N894, N649_0);
notg NOT1_156 (N895, N652_0);
notg NOT1_157 (N896, N655_0);
and_n #(2,0,0) AND2_158 (N897, {N49_1, N612_0});
and_n #(2,0,0) AND2_159 (N898, {N56_1, N608_0});
nand_n #(2,0,0) NAND2_160 (N899, {N53_1, N612_1});
nand_n #(2,0,0) NAND2_161 (N903, {N60_1, N608_1});
nand_n #(2,0,0) NAND2_162 (N907, {N49_2, N612_2});
nand_n #(2,0,0) NAND2_163 (N910, {N56_2, N608_2});
notg NOT1_164 (N913, N661_0);
notg NOT1_165 (N914, N658_0);
notg NOT1_166 (N915, N667_0);
notg NOT1_167 (N916, N664_0);
notg NOT1_168 (N917, N673_0);
notg NOT1_169 (N918, N670_0);
notg NOT1_170 (N919, N679_0);
notg NOT1_171 (N920, N676_0);
nand_n #(4,0,0) NAND4_172 (N921, {N277_1, N297_0, N326_2, N603_0});
nand_n #(4,0,0) NAND4_173 (N922, {N280_1, N297_1, N326_3, N603_1});
nand_n #(3,0,0) NAND3_174 (N923, {N303_0, N338_0, N603_2});
and_n #(3,0,0) AND3_175 (N926, {N303_1, N338_1, N603_3});
bufg BUFF1_176 (N935, N556_0);
notg NOT1_177 (N938, N688_0);
bufg BUFF1_178 (N939, N556_1);
notg NOT1_179 (N942, N691_0);
bufg BUFF1_180 (N943, N562_0);
notg NOT1_181 (N946, N694_0);
bufg BUFF1_182 (N947, N562_1);
notg NOT1_183 (N950, N697_0);
bufg BUFF1_184 (N951, N568_0);
notg NOT1_185 (N954, N700_0);
bufg BUFF1_186 (N955, N568_1);
notg NOT1_187 (N958, N703_0);
bufg BUFF1_188 (N959, N574_0);
bufg BUFF1_189 (N962, N574_1);
bufg BUFF1_190 (N965, N580_0);
notg NOT1_191 (N968, N706_0);
bufg BUFF1_192 (N969, N580_1);
notg NOT1_193 (N972, N709_0);
bufg BUFF1_194 (N973, N586_0);
notg NOT1_195 (N976, N712_0);
bufg BUFF1_196 (N977, N586_1);
notg NOT1_197 (N980, N715_0);
bufg BUFF1_198 (N981, N592_0);
notg NOT1_199 (N984, N628_0);
bufg BUFF1_200 (N985, N592_1);
notg NOT1_201 (N988, N718_0);
notg NOT1_202 (N989, N721_0);
notg NOT1_203 (N990, N634_0);
notg NOT1_204 (N991, N724_0);
notg NOT1_205 (N992, N727_0);
notg NOT1_206 (N993, N637_0);
bufg BUFF1_207 (N994, N595_0);
notg NOT1_208 (N997, N730_0);
bufg BUFF1_209 (N998, N595_1);
notg NOT1_210 (N1001, N733_0);
notg NOT1_211 (N1002, N736_0);
notg NOT1_212 (N1003, N739_0);
notg NOT1_213 (N1004, N640_0);
notg NOT1_214 (N1005, N742_0);
notg NOT1_215 (N1006, N745_0);
notg NOT1_216 (N1007, N646_0);
notg NOT1_217 (N1008, N748_0);
notg NOT1_218 (N1009, N751_0);
bufg BUFF1_219 (N1010, N559_0);
bufg BUFF1_220 (N1013, N559_1);
bufg BUFF1_221 (N1016, N565_0);
bufg BUFF1_222 (N1019, N565_1);
bufg BUFF1_223 (N1022, N571_0);
bufg BUFF1_224 (N1025, N571_1);
bufg BUFF1_225 (N1028, N577_0);
bufg BUFF1_226 (N1031, N577_1);
bufg BUFF1_227 (N1034, N583_0);
bufg BUFF1_228 (N1037, N583_1);
bufg BUFF1_229 (N1040, N589_0);
bufg BUFF1_230 (N1043, N589_1);
bufg BUFF1_231 (N1046, N598_0);
bufg BUFF1_232 (N1049, N598_1);
nand_n #(2,0,0) NAND2_233 (N1054, {N619_1, N888});
nand_n #(2,0,0) NAND2_234 (N1055, {N616_1, N889});
nand_n #(2,0,0) NAND2_235 (N1063, {N625_1, N890});
nand_n #(2,0,0) NAND2_236 (N1064, {N622_1, N891});
nand_n #(2,0,0) NAND2_237 (N1067, {N655_1, N895});
nand_n #(2,0,0) NAND2_238 (N1068, {N652_1, N896});
nand_n #(2,0,0) NAND2_239 (N1119, {N721_1, N988});
nand_n #(2,0,0) NAND2_240 (N1120, {N718_1, N989});
nand_n #(2,0,0) NAND2_241 (N1121, {N727_1, N991});
nand_n #(2,0,0) NAND2_242 (N1122, {N724_1, N992});
nand_n #(2,0,0) NAND2_243 (N1128, {N739_1, N1002});
nand_n #(2,0,0) NAND2_244 (N1129, {N736_1, N1003});
nand_n #(2,0,0) NAND2_245 (N1130, {N745_1, N1005});
nand_n #(2,0,0) NAND2_246 (N1131, {N742_1, N1006});
nand_n #(2,0,0) NAND2_247 (N1132, {N751_1, N1008});
nand_n #(2,0,0) NAND2_248 (N1133, {N748_1, N1009});
notg NOT1_249 (N1148, N939_0);
notg NOT1_250 (N1149, N935_0);
nand_n #(2,0,0) NAND2_251 (N1150, {N1054, N1055});
notg NOT1_252 (N1151, N943_0);
notg NOT1_253 (N1152, N947_0);
notg NOT1_254 (N1153, N955_0);
notg NOT1_255 (N1154, N951_0);
notg NOT1_256 (N1155, N962_0);
notg NOT1_257 (N1156, N969_0);
notg NOT1_258 (N1157, N977_0);
nand_n #(2,0,0) NAND2_259 (N1158, {N1063, N1064});
notg NOT1_260 (N1159, N985_0);
nand_n #(2,0,0) NAND2_261 (N1160, {N985_1, N892});
notg NOT1_262 (N1161, N998_0);
nand_n #(2,0,0) NAND2_263 (N1162, {N1067, N1068});
notg NOT1_264 (N1163, N899_0);
bufg BUFF1_265 (N1164, N899_1);
notg NOT1_266 (N1167, N903_0);
bufg BUFF1_267 (N1168, N903_1);
nand_n #(2,0,0) NAND2_268 (N1171, {N921, N923_0});
nand_n #(2,0,0) NAND2_269 (N1188, {N922, N923_1});
notg NOT1_270 (N1205, N1010_0);
nand_n #(2,0,0) NAND2_271 (N1206, {N1010_1, N938});
notg NOT1_272 (N1207, N1013_0);
nand_n #(2,0,0) NAND2_273 (N1208, {N1013_1, N942});
notg NOT1_274 (N1209, N1016_0);
nand_n #(2,0,0) NAND2_275 (N1210, {N1016_1, N946});
notg NOT1_276 (N1211, N1019_0);
nand_n #(2,0,0) NAND2_277 (N1212, {N1019_1, N950});
notg NOT1_278 (N1213, N1022_0);
nand_n #(2,0,0) NAND2_279 (N1214, {N1022_1, N954});
notg NOT1_280 (N1215, N1025_0);
nand_n #(2,0,0) NAND2_281 (N1216, {N1025_1, N958});
notg NOT1_282 (N1217, N1028_0);
notg NOT1_283 (N1218, N959_0);
notg NOT1_284 (N1219, N1031_0);
notg NOT1_285 (N1220, N1034_0);
nand_n #(2,0,0) NAND2_286 (N1221, {N1034_1, N968});
notg NOT1_287 (N1222, N965_0);
notg NOT1_288 (N1223, N1037_0);
nand_n #(2,0,0) NAND2_289 (N1224, {N1037_1, N972});
notg NOT1_290 (N1225, N1040_0);
nand_n #(2,0,0) NAND2_291 (N1226, {N1040_1, N976});
notg NOT1_292 (N1227, N973_0);
notg NOT1_293 (N1228, N1043_0);
nand_n #(2,0,0) NAND2_294 (N1229, {N1043_1, N980});
notg NOT1_295 (N1230, N981_0);
nand_n #(2,0,0) NAND2_296 (N1231, {N981_1, N984});
nand_n #(2,0,0) NAND2_297 (N1232, {N1119, N1120});
nand_n #(2,0,0) NAND2_298 (N1235, {N1121, N1122});
notg NOT1_299 (N1238, N1046_0);
nand_n #(2,0,0) NAND2_300 (N1239, {N1046_1, N997});
notg NOT1_301 (N1240, N994_0);
notg NOT1_302 (N1241, N1049_0);
nand_n #(2,0,0) NAND2_303 (N1242, {N1049_1, N1001});
nand_n #(2,0,0) NAND2_304 (N1243, {N1128, N1129});
nand_n #(2,0,0) NAND2_305 (N1246, {N1130, N1131});
nand_n #(2,0,0) NAND2_306 (N1249, {N1132, N1133});
bufg BUFF1_307 (N1252, N907_0);
bufg BUFF1_308 (N1255, N907_1);
bufg BUFF1_309 (N1258, N910_0);
bufg BUFF1_310 (N1261, N910_1);
notg NOT1_311 (N1264, N1150);
nand_n #(2,0,0) NAND2_312 (N1267, {N631_1, N1159});
nand_n #(2,0,0) NAND2_313 (N1309, {N688_1, N1205});
nand_n #(2,0,0) NAND2_314 (N1310, {N691_1, N1207});
nand_n #(2,0,0) NAND2_315 (N1311, {N694_1, N1209});
nand_n #(2,0,0) NAND2_316 (N1312, {N697_1, N1211});
nand_n #(2,0,0) NAND2_317 (N1313, {N700_1, N1213});
nand_n #(2,0,0) NAND2_318 (N1314, {N703_1, N1215});
nand_n #(2,0,0) NAND2_319 (N1315, {N706_1, N1220});
nand_n #(2,0,0) NAND2_320 (N1316, {N709_1, N1223});
nand_n #(2,0,0) NAND2_321 (N1317, {N712_1, N1225});
nand_n #(2,0,0) NAND2_322 (N1318, {N715_1, N1228});
notg NOT1_323 (N1319, N1158);
nand_n #(2,0,0) NAND2_324 (N1322, {N628_1, N1230});
nand_n #(2,0,0) NAND2_325 (N1327, {N730_1, N1238});
nand_n #(2,0,0) NAND2_326 (N1328, {N733_1, N1241});
notg NOT1_327 (N1334, N1162);
nand_n #(2,0,0) NAND2_328 (N1344, {N1267, N1160});
nand_n #(2,0,0) NAND2_329 (N1345, {N1249_0, N894});
notg NOT1_330 (N1346, N1249_1);
notg NOT1_331 (N1348, N1255_0);
notg NOT1_332 (N1349, N1252_0);
notg NOT1_333 (N1350, N1261_0);
notg NOT1_334 (N1351, N1258_0);
nand_n #(2,0,0) NAND2_335 (N1352, {N1309, N1206});
nand_n #(2,0,0) NAND2_336 (N1355, {N1310, N1208});
nand_n #(2,0,0) NAND2_337 (N1358, {N1311, N1210});
nand_n #(2,0,0) NAND2_338 (N1361, {N1312, N1212});
nand_n #(2,0,0) NAND2_339 (N1364, {N1313, N1214});
nand_n #(2,0,0) NAND2_340 (N1367, {N1314, N1216});
nand_n #(2,0,0) NAND2_341 (N1370, {N1315, N1221});
nand_n #(2,0,0) NAND2_342 (N1373, {N1316, N1224});
nand_n #(2,0,0) NAND2_343 (N1376, {N1317, N1226});
nand_n #(2,0,0) NAND2_344 (N1379, {N1318, N1229});
nand_n #(2,0,0) NAND2_345 (N1383, {N1322, N1231});
notg NOT1_346 (N1386, N1232_0);
nand_n #(2,0,0) NAND2_347 (N1387, {N1232_1, N990});
notg NOT1_348 (N1388, N1235_0);
nand_n #(2,0,0) NAND2_349 (N1389, {N1235_1, N993});
nand_n #(2,0,0) NAND2_350 (N1390, {N1327, N1239});
nand_n #(2,0,0) NAND2_351 (N1393, {N1328, N1242});
notg NOT1_352 (N1396, N1243_0);
nand_n #(2,0,0) NAND2_353 (N1397, {N1243_1, N1004});
notg NOT1_354 (N1398, N1246_0);
nand_n #(2,0,0) NAND2_355 (N1399, {N1246_1, N1007});
notg NOT1_356 (N1409, N1319_0);
nand_n #(2,0,0) NAND2_357 (N1412, {N649_1, N1346});
notg NOT1_358 (N1413, N1334_0);
bufg BUFF1_359 (N1416, N1264_0);
bufg BUFF1_360 (N1419, N1264_1);
nand_n #(2,0,0) NAND2_361 (N1433, {N634_1, N1386});
nand_n #(2,0,0) NAND2_362 (N1434, {N637_1, N1388});
nand_n #(2,0,0) NAND2_363 (N1438, {N640_1, N1396});
nand_n #(2,0,0) NAND2_364 (N1439, {N646_1, N1398});
notg NOT1_365 (N1440, N1344);
nand_n #(2,0,0) NAND2_366 (N1443, {N1355_0, N1148});
notg NOT1_367 (N1444, N1355_1);
nand_n #(2,0,0) NAND2_368 (N1445, {N1352_0, N1149});
notg NOT1_369 (N1446, N1352_1);
nand_n #(2,0,0) NAND2_370 (N1447, {N1358_0, N1151});
notg NOT1_371 (N1448, N1358_1);
nand_n #(2,0,0) NAND2_372 (N1451, {N1361_0, N1152});
notg NOT1_373 (N1452, N1361_1);
nand_n #(2,0,0) NAND2_374 (N1453, {N1367_0, N1153});
notg NOT1_375 (N1454, N1367_1);
nand_n #(2,0,0) NAND2_376 (N1455, {N1364_0, N1154});
notg NOT1_377 (N1456, N1364_1);
nand_n #(2,0,0) NAND2_378 (N1457, {N1373_0, N1156});
notg NOT1_379 (N1458, N1373_1);
nand_n #(2,0,0) NAND2_380 (N1459, {N1379_0, N1157});
notg NOT1_381 (N1460, N1379_1);
notg NOT1_382 (N1461, N1383_0);
nand_n #(2,0,0) NAND2_383 (N1462, {N1393_0, N1161});
notg NOT1_384 (N1463, N1393_1);
nand_n #(2,0,0) NAND2_385 (N1464, {N1345, N1412});
notg NOT1_386 (N1468, N1370_0);
nand_n #(2,0,0) NAND2_387 (N1469, {N1370_1, N1222});
notg NOT1_388 (N1470, N1376_0);
nand_n #(2,0,0) NAND2_389 (N1471, {N1376_1, N1227});
nand_n #(2,0,0) NAND2_390 (N1472, {N1387, N1433});
notg NOT1_391 (N1475, N1390_0);
nand_n #(2,0,0) NAND2_392 (N1476, {N1390_1, N1240});
nand_n #(2,0,0) NAND2_393 (N1478, {N1389, N1434});
nand_n #(2,0,0) NAND2_394 (N1481, {N1399, N1439});
nand_n #(2,0,0) NAND2_395 (N1484, {N1397, N1438});
nand_n #(2,0,0) NAND2_396 (N1487, {N939_1, N1444});
nand_n #(2,0,0) NAND2_397 (N1488, {N935_1, N1446});
nand_n #(2,0,0) NAND2_398 (N1489, {N943_1, N1448});
notg NOT1_399 (N1490, N1419_0);
notg NOT1_400 (N1491, N1416_0);
nand_n #(2,0,0) NAND2_401 (N1492, {N947_1, N1452});
nand_n #(2,0,0) NAND2_402 (N1493, {N955_1, N1454});
nand_n #(2,0,0) NAND2_403 (N1494, {N951_1, N1456});
nand_n #(2,0,0) NAND2_404 (N1495, {N969_1, N1458});
nand_n #(2,0,0) NAND2_405 (N1496, {N977_1, N1460});
nand_n #(2,0,0) NAND2_406 (N1498, {N998_1, N1463});
notg NOT1_407 (N1499, N1440_0);
nand_n #(2,0,0) NAND2_408 (N1500, {N965_1, N1468});
nand_n #(2,0,0) NAND2_409 (N1501, {N973_1, N1470});
nand_n #(2,0,0) NAND2_410 (N1504, {N994_1, N1475});
notg NOT1_411 (N1510, N1464);
nand_n #(2,0,0) NAND2_412 (N1513, {N1443, N1487});
nand_n #(2,0,0) NAND2_413 (N1514, {N1445, N1488});
nand_n #(2,0,0) NAND2_414 (N1517, {N1447, N1489});
nand_n #(2,0,0) NAND2_415 (N1520, {N1451, N1492});
nand_n #(2,0,0) NAND2_416 (N1521, {N1453, N1493});
nand_n #(2,0,0) NAND2_417 (N1522, {N1455, N1494});
nand_n #(2,0,0) NAND2_418 (N1526, {N1457, N1495});
nand_n #(2,0,0) NAND2_419 (N1527, {N1459, N1496});
notg NOT1_420 (N1528, N1472_0);
nand_n #(2,0,0) NAND2_421 (N1529, {N1462, N1498});
notg NOT1_422 (N1530, N1478_0);
notg NOT1_423 (N1531, N1481_0);
notg NOT1_424 (N1532, N1484_0);
nand_n #(2,0,0) NAND2_425 (N1534, {N1471, N1501});
nand_n #(2,0,0) NAND2_426 (N1537, {N1469, N1500});
nand_n #(2,0,0) NAND2_427 (N1540, {N1476, N1504});
notg NOT1_428 (N1546, N1513);
notg NOT1_429 (N1554, N1521);
notg NOT1_430 (N1557, N1526);
notg NOT1_431 (N1561, N1520);
nand_n #(2,0,0) NAND2_432 (N1567, {N1484_1, N1531});
nand_n #(2,0,0) NAND2_433 (N1568, {N1481_1, N1532});
notg NOT1_434 (N1569, N1510_0);
notg NOT1_435 (N1571, N1527);
notg NOT1_436 (N1576, N1529);
bufg BUFF1_437 (N1588, N1522_0);
notg NOT1_438 (N1591, N1534_0);
notg NOT1_439 (N1593, N1537_0);
nand_n #(2,0,0) NAND2_440 (N1594, {N1540_0, N1530});
notg NOT1_441 (N1595, N1540_1);
nand_n #(2,0,0) NAND2_442 (N1596, {N1567, N1568});
bufg BUFF1_443 (N1600, N1517_0);
bufg BUFF1_444 (N1603, N1517_1);
bufg BUFF1_445 (N1606, N1522_1);
bufg BUFF1_446 (N1609, N1522_2);
bufg BUFF1_447 (N1612, N1514_0);
bufg BUFF1_448 (N1615, N1514_1);
bufg BUFF1_449 (N1620, N1557_0);
bufg BUFF1_450 (N1623, N1554_0);
notg NOT1_451 (N1635, N1571_0);
nand_n #(2,0,0) NAND2_452 (N1636, {N1478_1, N1595});
nand_n #(2,0,0) NAND2_453 (N1638, {N1576_0, N1569});
notg NOT1_454 (N1639, N1576_1);
bufg BUFF1_455 (N1640, N1561_0);
bufg BUFF1_456 (N1643, N1561_1);
bufg BUFF1_457 (N1647, N1546_0);
bufg BUFF1_458 (N1651, N1546_1);
bufg BUFF1_459 (N1658, N1554_1);
bufg BUFF1_460 (N1661, N1557_1);
bufg BUFF1_461 (N1664, N1557_2);
nand_n #(2,0,0) NAND2_462 (N1671, {N1596_0, N893});
notg NOT1_463 (N1672, N1596_1);
notg NOT1_464 (N1675, N1600_0);
notg NOT1_465 (N1677, N1603_0);
nand_n #(2,0,0) NAND2_466 (N1678, {N1606_0, N1217});
notg NOT1_467 (N1679, N1606_1);
nand_n #(2,0,0) NAND2_468 (N1680, {N1609_0, N1219});
notg NOT1_469 (N1681, N1609_1);
notg NOT1_470 (N1682, N1612_0);
notg NOT1_471 (N1683, N1615_0);
nand_n #(2,0,0) NAND2_472 (N1685, {N1594, N1636});
nand_n #(2,0,0) NAND2_473 (N1688, {N1510_1, N1639});
bufg BUFF1_474 (N1697, N1588_0);
bufg BUFF1_475 (N1701, N1588_1);
nand_n #(2,0,0) NAND2_476 (N1706, {N643_1, N1672});
notg NOT1_477 (N1707, N1643_0);
nand_n #(2,0,0) NAND2_478 (N1708, {N1647_0, N1675});
notg NOT1_479 (N1709, N1647_1);
nand_n #(2,0,0) NAND2_480 (N1710, {N1651_0, N1677});
notg NOT1_481 (N1711, N1651_1);
nand_n #(2,0,0) NAND2_482 (N1712, {N1028_1, N1679});
nand_n #(2,0,0) NAND2_483 (N1713, {N1031_1, N1681});
bufg BUFF1_484 (N1714, N1620_0);
bufg BUFF1_485 (N1717, N1620_1);
nand_n #(2,0,0) NAND2_486 (N1720, {N1658_0, N1593});
notg NOT1_487 (N1721, N1658_1);
nand_n #(2,0,0) NAND2_488 (N1723, {N1638, N1688});
notg NOT1_489 (N1727, N1661_0);
notg NOT1_490 (N1728, N1640_0);
notg NOT1_491 (N1730, N1664_0);
bufg BUFF1_492 (N1731, N1623_0);
bufg BUFF1_493 (N1734, N1623_1);
nand_n #(2,0,0) NAND2_494 (N1740, {N1685_0, N1528});
notg NOT1_495 (N1741, N1685_1);
nand_n #(2,0,0) NAND2_496 (N1742, {N1671, N1706});
nand_n #(2,0,0) NAND2_497 (N1746, {N1600_1, N1709});
nand_n #(2,0,0) NAND2_498 (N1747, {N1603_1, N1711});
nand_n #(2,0,0) NAND2_499 (N1748, {N1678, N1712});
nand_n #(2,0,0) NAND2_500 (N1751, {N1680, N1713});
nand_n #(2,0,0) NAND2_501 (N1759, {N1537_1, N1721});
notg NOT1_502 (N1761, N1697_0);
nand_n #(2,0,0) NAND2_503 (N1762, {N1697_1, N1727});
notg NOT1_504 (N1763, N1701_0);
nand_n #(2,0,0) NAND2_505 (N1764, {N1701_1, N1730});
notg NOT1_506 (N1768, N1717_0);
nand_n #(2,0,0) NAND2_507 (N1769, {N1472_1, N1741});
nand_n #(2,0,0) NAND2_508 (N1772, {N1723_0, N1413});
notg NOT1_509 (N1773, N1723_1);
nand_n #(2,0,0) NAND2_510 (N1774, {N1708, N1746});
nand_n #(2,0,0) NAND2_511 (N1777, {N1710, N1747});
notg NOT1_512 (N1783, N1731_0);
nand_n #(2,0,0) NAND2_513 (N1784, {N1731_1, N1682});
notg NOT1_514 (N1785, N1714_0);
notg NOT1_515 (N1786, N1734_0);
nand_n #(2,0,0) NAND2_516 (N1787, {N1734_1, N1683});
nand_n #(2,0,0) NAND2_517 (N1788, {N1720, N1759});
nand_n #(2,0,0) NAND2_518 (N1791, {N1661_1, N1761});
nand_n #(2,0,0) NAND2_519 (N1792, {N1664_1, N1763});
nand_n #(2,0,0) NAND2_520 (N1795, {N1751_0, N1155});
notg NOT1_521 (N1796, N1751_1);
nand_n #(2,0,0) NAND2_522 (N1798, {N1740, N1769});
nand_n #(2,0,0) NAND2_523 (N1801, {N1334_1, N1773});
nand_n #(2,0,0) NAND2_524 (N1802, {N1742_0, N290_0});
notg NOT1_525 (N1807, N1748_0);
nand_n #(2,0,0) NAND2_526 (N1808, {N1748_1, N1218});
nand_n #(2,0,0) NAND2_527 (N1809, {N1612_1, N1783});
nand_n #(2,0,0) NAND2_528 (N1810, {N1615_1, N1786});
nand_n #(2,0,0) NAND2_529 (N1812, {N1791, N1762});
nand_n #(2,0,0) NAND2_530 (N1815, {N1792, N1764});
bufg BUFF1_531 (N1818, N1742_1);
nand_n #(2,0,0) NAND2_532 (N1821, {N1777_0, N1490});
notg NOT1_533 (N1822, N1777_1);
nand_n #(2,0,0) NAND2_534 (N1823, {N1774_0, N1491});
notg NOT1_535 (N1824, N1774_1);
nand_n #(2,0,0) NAND2_536 (N1825, {N962_1, N1796});
nand_n #(2,0,0) NAND2_537 (N1826, {N1788_0, N1409});
notg NOT1_538 (N1827, N1788_1);
nand_n #(2,0,0) NAND2_539 (N1830, {N1772, N1801});
nand_n #(2,0,0) NAND2_540 (N1837, {N959_1, N1807});
nand_n #(2,0,0) NAND2_541 (N1838, {N1809, N1784});
nand_n #(2,0,0) NAND2_542 (N1841, {N1810, N1787});
nand_n #(2,0,0) NAND2_543 (N1848, {N1419_1, N1822});
nand_n #(2,0,0) NAND2_544 (N1849, {N1416_1, N1824});
nand_n #(2,0,0) NAND2_545 (N1850, {N1795, N1825});
nand_n #(2,0,0) NAND2_546 (N1852, {N1319_1, N1827});
nand_n #(2,0,0) NAND2_547 (N1855, {N1815_0, N1707});
notg NOT1_548 (N1856, N1815_1);
notg NOT1_549 (N1857, N1818_0);
nand_n #(2,0,0) NAND2_550 (N1858, {N1798_0, N290_1});
notg NOT1_551 (N1864, N1812_0);
nand_n #(2,0,0) NAND2_552 (N1865, {N1812_1, N1728});
bufg BUFF1_553 (N1866, N1798_1);
bufg BUFF1_554 (N1869, N1802_0);
bufg BUFF1_555 (N1872, N1802_1);
nand_n #(2,0,0) NAND2_556 (N1875, {N1808, N1837});
nand_n #(2,0,0) NAND2_557 (N1878, {N1821, N1848});
nand_n #(2,0,0) NAND2_558 (N1879, {N1823, N1849});
nand_n #(2,0,0) NAND2_559 (N1882, {N1841_0, N1768});
notg NOT1_560 (N1883, N1841_1);
nand_n #(2,0,0) NAND2_561 (N1884, {N1826, N1852});
nand_n #(2,0,0) NAND2_562 (N1885, {N1643_1, N1856});
nand_n #(2,0,0) NAND2_563 (N1889, {N1830_0, N290_2});
notg NOT1_564 (N1895, N1838_0);
nand_n #(2,0,0) NAND2_565 (N1896, {N1838_1, N1785});
nand_n #(2,0,0) NAND2_566 (N1897, {N1640_1, N1864});
notg NOT1_567 (N1898, N1850);
bufg BUFF1_568 (N1902, N1830_1);
notg NOT1_569 (N1910, N1878);
nand_n #(2,0,0) NAND2_570 (N1911, {N1717_1, N1883});
notg NOT1_571 (N1912, N1884);
nand_n #(2,0,0) NAND2_572 (N1913, {N1855, N1885});
notg NOT1_573 (N1915, N1866_0);
nand_n #(2,0,0) NAND2_574 (N1919, {N1872_0, N919});
notg NOT1_575 (N1920, N1872_1);
nand_n #(2,0,0) NAND2_576 (N1921, {N1869_0, N920});
notg NOT1_577 (N1922, N1869_1);
notg NOT1_578 (N1923, N1875_0);
nand_n #(2,0,0) NAND2_579 (N1924, {N1714_1, N1895});
bufg BUFF1_580 (N1927, N1858_0);
bufg BUFF1_581 (N1930, N1858_1);
nand_n #(2,0,0) NAND2_582 (N1933, {N1865, N1897});
nand_n #(2,0,0) NAND2_583 (N1936, {N1882, N1911});
notg NOT1_584 (N1937, N1898_0);
notg NOT1_585 (N1938, N1902_0);
nand_n #(2,0,0) NAND2_586 (N1941, {N679_1, N1920});
nand_n #(2,0,0) NAND2_587 (N1942, {N676_1, N1922});
bufg BUFF1_588 (N1944, N1879_0);
notg NOT1_589 (N1947, N1913);
bufg BUFF1_590 (N1950, N1889_0);
bufg BUFF1_591 (N1953, N1889_1);
bufg BUFF1_592 (N1958, N1879_1);
nand_n #(2,0,0) NAND2_593 (N1961, {N1896, N1924});
and_n #(2,0,0) AND2_594 (N1965, {N1910, N601});
and_n #(2,0,0) AND2_595 (N1968, {N602, N1912});
nand_n #(2,0,0) NAND2_596 (N1975, {N1930_0, N917});
notg NOT1_597 (N1976, N1930_1);
nand_n #(2,0,0) NAND2_598 (N1977, {N1927_0, N918});
notg NOT1_599 (N1978, N1927_1);
nand_n #(2,0,0) NAND2_600 (N1979, {N1919, N1941});
nand_n #(2,0,0) NAND2_601 (N1980, {N1921, N1942});
notg NOT1_602 (N1985, N1933_0);
notg NOT1_603 (N1987, N1936);
notg NOT1_604 (N1999, N1944_0);
nand_n #(2,0,0) NAND2_605 (N2000, {N1944_1, N1937});
notg NOT1_606 (N2002, N1947_0);
nand_n #(2,0,0) NAND2_607 (N2003, {N1947_1, N1499});
nand_n #(2,0,0) NAND2_608 (N2004, {N1953_0, N1350});
notg NOT1_609 (N2005, N1953_1);
nand_n #(2,0,0) NAND2_610 (N2006, {N1950_0, N1351});
notg NOT1_611 (N2007, N1950_1);
nand_n #(2,0,0) NAND2_612 (N2008, {N673_1, N1976});
nand_n #(2,0,0) NAND2_613 (N2009, {N670_1, N1978});
notg NOT1_614 (N2012, N1979);
notg NOT1_615 (N2013, N1958_0);
nand_n #(2,0,0) NAND2_616 (N2014, {N1958_1, N1923});
notg NOT1_617 (N2015, N1961_0);
nand_n #(2,0,0) NAND2_618 (N2016, {N1961_1, N1635});
notg NOT1_619 (N2018, N1965_0);
notg NOT1_620 (N2019, N1968_0);
nand_n #(2,0,0) NAND2_621 (N2020, {N1898_1, N1999});
notg NOT1_622 (N2021, N1987_0);
nand_n #(2,0,0) NAND2_623 (N2022, {N1987_1, N1591});
nand_n #(2,0,0) NAND2_624 (N2023, {N1440_1, N2002});
nand_n #(2,0,0) NAND2_625 (N2024, {N1261_1, N2005});
nand_n #(2,0,0) NAND2_626 (N2025, {N1258_1, N2007});
nand_n #(2,0,0) NAND2_627 (N2026, {N1975, N2008});
nand_n #(2,0,0) NAND2_628 (N2027, {N1977, N2009});
notg NOT1_629 (N2030, N1980_0);
bufg BUFF1_630 (N2033, N1980_1);
nand_n #(2,0,0) NAND2_631 (N2036, {N1875_1, N2013});
nand_n #(2,0,0) NAND2_632 (N2037, {N1571_1, N2015});
nand_n #(2,0,0) NAND2_633 (N2038, {N2020, N2000});
nand_n #(2,0,0) NAND2_634 (N2039, {N1534_1, N2021});
nand_n #(2,0,0) NAND2_635 (N2040, {N2023, N2003});
nand_n #(2,0,0) NAND2_636 (N2041, {N2004, N2024});
nand_n #(2,0,0) NAND2_637 (N2042, {N2006, N2025});
notg NOT1_638 (N2047, N2026);
nand_n #(2,0,0) NAND2_639 (N2052, {N2036, N2014});
nand_n #(2,0,0) NAND2_640 (N2055, {N2037, N2016});
notg NOT1_641 (N2060, N2038);
nand_n #(2,0,0) NAND2_642 (N2061, {N2039, N2022});
nand_n #(2,0,0) NAND2_643 (N2062, {N2040, N290_3});
notg NOT1_644 (N2067, N2041);
notg NOT1_645 (N2068, N2027_0);
bufg BUFF1_646 (N2071, N2027_1);
notg NOT1_647 (N2076, N2052_0);
notg NOT1_648 (N2077, N2055_0);
nand_n #(2,0,0) NAND2_649 (N2078, {N2060, N290_4});
nand_n #(2,0,0) NAND2_650 (N2081, {N2061, N290_5});
notg NOT1_651 (N2086, N2042_0);
bufg BUFF1_652 (N2089, N2042_1);
and_n #(2,0,0) AND2_653 (N2104, {N2030_0, N2068_0});
and_n #(2,0,0) AND2_654 (N2119, {N2033_0, N2068_1});
and_n #(2,0,0) AND2_655 (N2129, {N2030_1, N2071_0});
and_n #(2,0,0) AND2_656 (N2143, {N2033_1, N2071_1});
bufg BUFF1_657 (N2148, N2062_0);
bufg BUFF1_658 (N2151, N2062_1);
bufg BUFF1_659 (N2196, N2078_0);
bufg BUFF1_660 (N2199, N2078_1);
bufg BUFF1_661 (N2202, N2081_0);
bufg BUFF1_662 (N2205, N2081_1);
nand_n #(2,0,0) NAND2_663 (N2214, {N2151_0, N915});
notg NOT1_664 (N2215, N2151_1);
nand_n #(2,0,0) NAND2_665 (N2216, {N2148_0, N916});
notg NOT1_666 (N2217, N2148_1);
nand_n #(2,0,0) NAND2_667 (N2222, {N2199_0, N1348});
notg NOT1_668 (N2223, N2199_1);
nand_n #(2,0,0) NAND2_669 (N2224, {N2196_0, N1349});
notg NOT1_670 (N2225, N2196_1);
nand_n #(2,0,0) NAND2_671 (N2226, {N2205_0, N913});
notg NOT1_672 (N2227, N2205_1);
nand_n #(2,0,0) NAND2_673 (N2228, {N2202_0, N914});
notg NOT1_674 (N2229, N2202_1);
nand_n #(2,0,0) NAND2_675 (N2230, {N667_1, N2215});
nand_n #(2,0,0) NAND2_676 (N2231, {N664_1, N2217});
nand_n #(2,0,0) NAND2_677 (N2232, {N1255_1, N2223});
nand_n #(2,0,0) NAND2_678 (N2233, {N1252_1, N2225});
nand_n #(2,0,0) NAND2_679 (N2234, {N661_1, N2227});
nand_n #(2,0,0) NAND2_680 (N2235, {N658_1, N2229});
nand_n #(2,0,0) NAND2_681 (N2236, {N2214, N2230});
nand_n #(2,0,0) NAND2_682 (N2237, {N2216, N2231});
nand_n #(2,0,0) NAND2_683 (N2240, {N2222, N2232});
nand_n #(2,0,0) NAND2_684 (N2241, {N2224, N2233});
nand_n #(2,0,0) NAND2_685 (N2244, {N2226, N2234});
nand_n #(2,0,0) NAND2_686 (N2245, {N2228, N2235});
notg NOT1_687 (N2250, N2236);
notg NOT1_688 (N2253, N2240);
notg NOT1_689 (N2256, N2244);
notg NOT1_690 (N2257, N2237_0);
bufg BUFF1_691 (N2260, N2237_1);
notg NOT1_692 (N2263, N2241_0);
and_n #(2,0,0) AND2_693 (N2266, {N1164_0, N2241_1});
notg NOT1_694 (N2269, N2245_0);
and_n #(2,0,0) AND2_695 (N2272, {N1168_0, N2245_1});
nand_n #(8,0,0) NAND8_696 (N2279, {N2067, N2012, N2047, N2250, N899_2, N2256, N2253, N903_2});
bufg BUFF1_697 (N2286, N2266_0);
bufg BUFF1_698 (N2297, N2266_1);
bufg BUFF1_699 (N2315, N2272_0);
bufg BUFF1_700 (N2326, N2272_1);
and_n #(2,0,0) AND2_701 (N2340, {N2086_0, N2257_0});
and_n #(2,0,0) AND2_702 (N2353, {N2089_0, N2257_1});
and_n #(2,0,0) AND2_703 (N2361, {N2086_1, N2260_0});
and_n #(2,0,0) AND2_704 (N2375, {N2089_1, N2260_1});
and_n #(4,0,0) AND4_705 (N2384, {N338_2, N2279_0, N313_0, N313_1});
and_n #(2,0,0) AND2_706 (N2385, {N1163, N2263_0});
and_n #(2,0,0) AND2_707 (N2386, {N1164_1, N2263_1});
and_n #(2,0,0) AND2_708 (N2426, {N1167, N2269_0});
and_n #(2,0,0) AND2_709 (N2427, {N1168_1, N2269_1});
nand_n #(5,0,0) NAND5_710 (N2537, {N2286_0, N2315_0, N2361_0, N2104_0, N1171_0});
nand_n #(5,0,0) NAND5_711 (N2540, {N2286_1, N2315_1, N2340_0, N2129_0, N1171_1});
nand_n #(5,0,0) NAND5_712 (N2543, {N2286_2, N2315_2, N2340_1, N2119_0, N1171_2});
nand_n #(5,0,0) NAND5_713 (N2546, {N2286_3, N2315_3, N2353_0, N2104_1, N1171_3});
nand_n #(5,0,0) NAND5_714 (N2549, {N2297_0, N2315_4, N2375_0, N2119_1, N1188_0});
nand_n #(5,0,0) NAND5_715 (N2552, {N2297_1, N2326_0, N2361_1, N2143_0, N1188_1});
nand_n #(5,0,0) NAND5_716 (N2555, {N2297_2, N2326_1, N2375_1, N2129_1, N1188_2});
and_n #(5,0,0) AND5_717 (N2558, {N2286_4, N2315_5, N2361_2, N2104_2, N1171_4});
and_n #(5,0,0) AND5_718 (N2561, {N2286_5, N2315_6, N2340_2, N2129_2, N1171_5});
and_n #(5,0,0) AND5_719 (N2564, {N2286_6, N2315_7, N2340_3, N2119_2, N1171_6});
and_n #(5,0,0) AND5_720 (N2567, {N2286_7, N2315_8, N2353_1, N2104_3, N1171_7});
and_n #(5,0,0) AND5_721 (N2570, {N2297_3, N2315_9, N2375_2, N2119_3, N1188_3});
and_n #(5,0,0) AND5_722 (N2573, {N2297_4, N2326_2, N2361_3, N2143_1, N1188_4});
and_n #(5,0,0) AND5_723 (N2576, {N2297_5, N2326_3, N2375_3, N2129_3, N1188_5});
nand_n #(5,0,0) NAND5_724 (N2594, {N2286_8, N2427_0, N2361_4, N2129_4, N1171_8});
nand_n #(5,0,0) NAND5_725 (N2597, {N2297_6, N2427_1, N2361_5, N2119_4, N1171_9});
nand_n #(5,0,0) NAND5_726 (N2600, {N2297_7, N2427_2, N2375_4, N2104_4, N1171_10});
nand_n #(5,0,0) NAND5_727 (N2603, {N2297_8, N2427_3, N2340_4, N2143_2, N1171_11});
nand_n #(5,0,0) NAND5_728 (N2606, {N2297_9, N2427_4, N2353_2, N2129_5, N1188_6});
nand_n #(5,0,0) NAND5_729 (N2611, {N2386_0, N2326_4, N2361_6, N2129_6, N1188_7});
nand_n #(5,0,0) NAND5_730 (N2614, {N2386_1, N2326_5, N2361_7, N2119_5, N1188_8});
nand_n #(5,0,0) NAND5_731 (N2617, {N2386_2, N2326_6, N2375_5, N2104_5, N1188_9});
nand_n #(5,0,0) NAND5_732 (N2620, {N2386_3, N2326_7, N2353_3, N2129_7, N1188_10});
nand_n #(5,0,0) NAND5_733 (N2627, {N2297_10, N2427_5, N2340_5, N2104_6, N926_0});
nand_n #(5,0,0) NAND5_734 (N2628, {N2386_4, N2326_8, N2340_6, N2104_7, N926_1});
nand_n #(5,0,0) NAND5_735 (N2629, {N2386_5, N2427_6, N2361_8, N2104_8, N926_2});
nand_n #(5,0,0) NAND5_736 (N2630, {N2386_6, N2427_7, N2340_7, N2129_8, N926_3});
nand_n #(5,0,0) NAND5_737 (N2631, {N2386_7, N2427_8, N2340_8, N2119_6, N926_4});
nand_n #(5,0,0) NAND5_738 (N2632, {N2386_8, N2427_9, N2353_4, N2104_9, N926_5});
nand_n #(5,0,0) NAND5_739 (N2633, {N2386_9, N2426, N2340_9, N2104_10, N926_6});
nand_n #(5,0,0) NAND5_740 (N2634, {N2385, N2427_10, N2340_10, N2104_11, N926_7});
and_n #(5,0,0) AND5_741 (N2639, {N2286_9, N2427_11, N2361_9, N2129_9, N1171_12});
and_n #(5,0,0) AND5_742 (N2642, {N2297_11, N2427_12, N2361_10, N2119_7, N1171_13});
and_n #(5,0,0) AND5_743 (N2645, {N2297_12, N2427_13, N2375_6, N2104_12, N1171_14});
and_n #(5,0,0) AND5_744 (N2648, {N2297_13, N2427_14, N2340_11, N2143_3, N1171_15});
and_n #(5,0,0) AND5_745 (N2651, {N2297_14, N2427_15, N2353_5, N2129_10, N1188_11});
and_n #(5,0,0) AND5_746 (N2655, {N2386_10, N2326_9, N2361_11, N2129_11, N1188_12});
and_n #(5,0,0) AND5_747 (N2658, {N2386_11, N2326_10, N2361_12, N2119_8, N1188_13});
and_n #(5,0,0) AND5_748 (N2661, {N2386_12, N2326_11, N2375_7, N2104_13, N1188_14});
and_n #(5,0,0) AND5_749 (N2664, {N2386_13, N2326_12, N2353_6, N2129_12, N1188_15});
nand_n #(2,0,0) NAND2_750 (N2669, {N2558_0, N534});
notg NOT1_751 (N2670, N2558_1);
nand_n #(2,0,0) NAND2_752 (N2671, {N2561_0, N535});
notg NOT1_753 (N2672, N2561_1);
nand_n #(2,0,0) NAND2_754 (N2673, {N2564_0, N536});
notg NOT1_755 (N2674, N2564_1);
nand_n #(2,0,0) NAND2_756 (N2675, {N2567_0, N537});
notg NOT1_757 (N2676, N2567_1);
nand_n #(2,0,0) NAND2_758 (N2682, {N2570_0, N543});
notg NOT1_759 (N2683, N2570_1);
nand_n #(2,0,0) NAND2_760 (N2688, {N2573_0, N548});
notg NOT1_761 (N2689, N2573_1);
nand_n #(2,0,0) NAND2_762 (N2690, {N2576_0, N549});
notg NOT1_763 (N2691, N2576_1);
and_n #(8,0,0) AND8_764 (N2710, {N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634});
nand_n #(2,0,0) NAND2_765 (N2720, {N343_1, N2670});
nand_n #(2,0,0) NAND2_766 (N2721, {N346_1, N2672});
nand_n #(2,0,0) NAND2_767 (N2722, {N349_1, N2674});
nand_n #(2,0,0) NAND2_768 (N2723, {N352_1, N2676});
nand_n #(2,0,0) NAND2_769 (N2724, {N2639_0, N538});
notg NOT1_770 (N2725, N2639_1);
nand_n #(2,0,0) NAND2_771 (N2726, {N2642_0, N539});
notg NOT1_772 (N2727, N2642_1);
nand_n #(2,0,0) NAND2_773 (N2728, {N2645_0, N540});
notg NOT1_774 (N2729, N2645_1);
nand_n #(2,0,0) NAND2_775 (N2730, {N2648_0, N541});
notg NOT1_776 (N2731, N2648_1);
nand_n #(2,0,0) NAND2_777 (N2732, {N2651_0, N542});
notg NOT1_778 (N2733, N2651_1);
nand_n #(2,0,0) NAND2_779 (N2734, {N370_1, N2683});
nand_n #(2,0,0) NAND2_780 (N2735, {N2655_0, N544});
notg NOT1_781 (N2736, N2655_1);
nand_n #(2,0,0) NAND2_782 (N2737, {N2658_0, N545});
notg NOT1_783 (N2738, N2658_1);
nand_n #(2,0,0) NAND2_784 (N2739, {N2661_0, N546});
notg NOT1_785 (N2740, N2661_1);
nand_n #(2,0,0) NAND2_786 (N2741, {N2664_0, N547});
notg NOT1_787 (N2742, N2664_1);
nand_n #(2,0,0) NAND2_788 (N2743, {N385_1, N2689});
nand_n #(2,0,0) NAND2_789 (N2744, {N388_1, N2691});
nand_n #(8,0,0) NAND8_790 (N2745, {N2537_0, N2540_0, N2543_0, N2546_0, N2594_0, N2597_0, N2600_0, N2603_0});
nand_n #(8,0,0) NAND8_791 (N2746, {N2606_0, N2549_0, N2611_0, N2614_0, N2617_0, N2620_0, N2552_0, N2555_0});
and_n #(8,0,0) AND8_792 (N2747, {N2537_1, N2540_1, N2543_1, N2546_1, N2594_1, N2597_1, N2600_1, N2603_1});
and_n #(8,0,0) AND8_793 (N2750, {N2606_1, N2549_1, N2611_1, N2614_1, N2617_1, N2620_1, N2552_1, N2555_1});
nand_n #(2,0,0) NAND2_794 (N2753, {N2669, N2720});
nand_n #(2,0,0) NAND2_795 (N2754, {N2671, N2721});
nand_n #(2,0,0) NAND2_796 (N2755, {N2673, N2722});
nand_n #(2,0,0) NAND2_797 (N2756, {N2675, N2723});
nand_n #(2,0,0) NAND2_798 (N2757, {N355_1, N2725});
nand_n #(2,0,0) NAND2_799 (N2758, {N358_1, N2727});
nand_n #(2,0,0) NAND2_800 (N2759, {N361_1, N2729});
nand_n #(2,0,0) NAND2_801 (N2760, {N364_1, N2731});
nand_n #(2,0,0) NAND2_802 (N2761, {N367_1, N2733});
nand_n #(2,0,0) NAND2_803 (N2762, {N2682, N2734});
nand_n #(2,0,0) NAND2_804 (N2763, {N373_1, N2736});
nand_n #(2,0,0) NAND2_805 (N2764, {N376_1, N2738});
nand_n #(2,0,0) NAND2_806 (N2765, {N379_1, N2740});
nand_n #(2,0,0) NAND2_807 (N2766, {N382_1, N2742});
nand_n #(2,0,0) NAND2_808 (N2767, {N2688, N2743});
nand_n #(2,0,0) NAND2_809 (N2768, {N2690, N2744});
and_n #(2,0,0) AND2_810 (N2773, {N2745, N275});
and_n #(2,0,0) AND2_811 (N2776, {N2746, N276});
nand_n #(2,0,0) NAND2_812 (N2779, {N2724, N2757});
nand_n #(2,0,0) NAND2_813 (N2780, {N2726, N2758});
nand_n #(2,0,0) NAND2_814 (N2781, {N2728, N2759});
nand_n #(2,0,0) NAND2_815 (N2782, {N2730, N2760});
nand_n #(2,0,0) NAND2_816 (N2783, {N2732, N2761});
nand_n #(2,0,0) NAND2_817 (N2784, {N2735, N2763});
nand_n #(2,0,0) NAND2_818 (N2785, {N2737, N2764});
nand_n #(2,0,0) NAND2_819 (N2786, {N2739, N2765});
nand_n #(2,0,0) NAND2_820 (N2787, {N2741, N2766});
and_n #(3,0,0) AND3_821 (N2788, {N2747_0, N2750_0, N2710});
nand_n #(2,0,0) NAND2_822 (N2789, {N2747_1, N2750_1});
and_n #(4,0,0) AND4_823 (N2800, {N338_3, N2279_1, N99_3, N2788});
nand_n #(2,0,0) NAND2_824 (N2807, {N2773_0, N2018});
notg NOT1_825 (N2808, N2773_1);
nand_n #(2,0,0) NAND2_826 (N2809, {N2776_0, N2019});
notg NOT1_827 (N2810, N2776_1);
nor_n #(2,0,0) NOR2_828 (N2811, {N2384, N2800});
and_n #(3,0,0) AND3_829 (N2812, {N897, N283_0, N2789_0});
and_n #(3,0,0) AND3_830 (N2815, {N76_1, N283_1, N2789_1});
and_n #(3,0,0) AND3_831 (N2818, {N82_1, N283_2, N2789_2});
and_n #(3,0,0) AND3_832 (N2821, {N85_1, N283_3, N2789_3});
and_n #(3,0,0) AND3_833 (N2824, {N898, N283_4, N2789_4});
nand_n #(2,0,0) NAND2_834 (N2827, {N1965_1, N2808});
nand_n #(2,0,0) NAND2_835 (N2828, {N1968_1, N2810});
and_n #(3,0,0) AND3_836 (N2829, {N79_1, N283_5, N2789_5});
nand_n #(2,0,0) NAND2_837 (N2843, {N2807, N2827});
nand_n #(2,0,0) NAND2_838 (N2846, {N2809, N2828});
nand_n #(2,0,0) NAND2_839 (N2850, {N2812_0, N2076});
nand_n #(2,0,0) NAND2_840 (N2851, {N2815_0, N2077});
nand_n #(2,0,0) NAND2_841 (N2852, {N2818_0, N1915});
nand_n #(2,0,0) NAND2_842 (N2853, {N2821_0, N1857});
nand_n #(2,0,0) NAND2_843 (N2854, {N2824_0, N1938});
notg NOT1_844 (N2857, N2812_1);
notg NOT1_845 (N2858, N2815_1);
notg NOT1_846 (N2859, N2818_1);
notg NOT1_847 (N2860, N2821_1);
notg NOT1_848 (N2861, N2824_1);
notg NOT1_849 (N2862, N2829_0);
nand_n #(2,0,0) NAND2_850 (N2863, {N2829_1, N1985});
nand_n #(2,0,0) NAND2_851 (N2866, {N2052_1, N2857});
nand_n #(2,0,0) NAND2_852 (N2867, {N2055_1, N2858});
nand_n #(2,0,0) NAND2_853 (N2868, {N1866_1, N2859});
nand_n #(2,0,0) NAND2_854 (N2869, {N1818_1, N2860});
nand_n #(2,0,0) NAND2_855 (N2870, {N1902_1, N2861});
nand_n #(2,0,0) NAND2_856 (N2871, {N2843_0, N886});
notg NOT1_857 (N2872, N2843_1);
nand_n #(2,0,0) NAND2_858 (N2873, {N2846_0, N887});
notg NOT1_859 (N2874, N2846_1);
nand_n #(2,0,0) NAND2_860 (N2875, {N1933_1, N2862});
nand_n #(2,0,0) NAND2_861 (N2876, {N2866, N2850});
nand_n #(2,0,0) NAND2_862 (N2877, {N2867, N2851});
nand_n #(2,0,0) NAND2_863 (N2878, {N2868, N2852});
nand_n #(2,0,0) NAND2_864 (N2879, {N2869, N2853});
nand_n #(2,0,0) NAND2_865 (N2880, {N2870, N2854});
nand_n #(2,0,0) NAND2_866 (N2881, {N682_1, N2872});
nand_n #(2,0,0) NAND2_867 (N2882, {N685_1, N2874});
nand_n #(2,0,0) NAND2_868 (N2883, {N2875, N2863});
and_n #(2,0,0) AND2_869 (N2886, {N2876, N550});
and_n #(2,0,0) AND2_870 (N2887, {N551, N2877});
and_n #(2,0,0) AND2_871 (N2888, {N553, N2878});
and_n #(2,0,0) AND2_872 (N2889, {N2879, N554});
and_n #(2,0,0) AND2_873 (N2890, {N555, N2880});
nand_n #(2,0,0) NAND2_874 (N2891, {N2871, N2881});
nand_n #(2,0,0) NAND2_875 (N2892, {N2873, N2882});
nand_n #(2,0,0) NAND2_876 (N2895, {N2883_0, N1461});
notg NOT1_877 (N2896, N2883_1);
nand_n #(2,0,0) NAND2_878 (N2897, {N1383_1, N2896});
nand_n #(2,0,0) NAND2_879 (N2898, {N2895, N2897});
and_n #(2,0,0) AND2_880 (N2899, {N2898, N552});

endmodule
