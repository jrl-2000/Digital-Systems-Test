/****************************************************************************
 *                                                                          *
 *  FLAT VERSION of HIGH-LEVEL MODEL for c3540                              *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *  Verified  by: Jonathan David Hauke (jhauke@eecs.umich.edu)              *
 *                                                                          *
 *                Oct 20, 1998                                              *
 *                                                                          *
****************************************************************************/

// Flat Verilog File 
module c3540g (
	in50, in58, in68, in77, in87, in97, in107, 
	in116, in226, in232, in238, in244, in250, in257, in264, 
	in270, in124, in125, in128, in132, in137, in143, in150, 
	in159, in283, in294, in303, in311, in317, in322, in326, 
	in329, in222, in223, in330, in274, in2897, in200, in190, 
	in179, in343, in213, in169, in45, in41, in1698, in33, 
	in20, in13, in1,
	out375, out378, out381, out384, out387, out390, out393, 
	out396, out407, out409, out402, out351, out358, out405, out399, 
	out369, out372, out353, out355, out361, out364, out367);

   input
	in50, in58, in68, in77, in87, in97, in107, 
	in116, in226, in232, in238, in244, in250, in257, in264, 
	in270, in124, in125, in128, in132, in137, in143, in150, 
	in159, in283, in294, in303, in311, in317, in322, in326, 
	in329, in222, in223, in330, in274, in2897, in200, in190, 
	in179, in343, in213, in169, in45, in41, in1698, in33, 
	in20, in13, in1;

   output
	out375, out378, out381, out384, out387, out390, out393, 
	out396, out407, out409, out402, out351, out358, out405, out399, 
	out369, out372, out353, out355, out361, out364, out367;

inv M1_UM1_0_BaD0(in107, A_BCDbus_1);
inv M1_UM1_0_BaD1_Xo0(in97, M1_UM1_0_BaD1_NotA);
inv M1_UM1_0_BaD1_Xo1(in107, M1_UM1_0_BaD1_NotB);
nand2 M1_UM1_0_BaD1_Xo2(M1_UM1_0_BaD1_NotA, in107, M1_UM1_0_BaD1_line2);
nand2 M1_UM1_0_BaD1_Xo3(M1_UM1_0_BaD1_NotB, in97, M1_UM1_0_BaD1_line3);
nand2 M1_UM1_0_BaD1_Xo4(M1_UM1_0_BaD1_line2, M1_UM1_0_BaD1_line3, M1_UM1_0_line1);
inv M1_UM1_0_BaD2(M1_UM1_0_line1, A_BCDbus_2);
inv M1_UM1_0_BaD3(in97, M1_UM1_0_line3);
inv M1_UM1_0_BaD4(in87, M1_UM1_0_line4);
nand3 M1_UM1_0_BaD5(A_BCDbus_1, M1_UM1_0_line3, M1_UM1_0_line4, A_BCDbus_3);
inv M1_UM1_1_BaD0(in68, A_BCDbus_5);
inv M1_UM1_1_BaD1_Xo0(in58, M1_UM1_1_BaD1_NotA);
inv M1_UM1_1_BaD1_Xo1(in68, M1_UM1_1_BaD1_NotB);
nand2 M1_UM1_1_BaD1_Xo2(M1_UM1_1_BaD1_NotA, in68, M1_UM1_1_BaD1_line2);
nand2 M1_UM1_1_BaD1_Xo3(M1_UM1_1_BaD1_NotB, in58, M1_UM1_1_BaD1_line3);
nand2 M1_UM1_1_BaD1_Xo4(M1_UM1_1_BaD1_line2, M1_UM1_1_BaD1_line3, M1_UM1_1_line1);
inv M1_UM1_1_BaD2(M1_UM1_1_line1, A_BCDbus_6);
inv M1_UM1_1_BaD3(in58, M1_UM1_1_line3);
inv M1_UM1_1_BaD4(in50, M1_UM1_1_line4);
nand3 M1_UM1_1_BaD5(A_BCDbus_5, M1_UM1_1_line3, M1_UM1_1_line4, A_BCDbus_7);
inv M2_Inv8_0_Inv4_0(in116, Not_Abus_0);
inv M2_Inv8_0_Inv4_1(in107, Not_Abus_1);
inv M2_Inv8_0_Inv4_2(in97, Not_Abus_2);
inv M2_Inv8_0_Inv4_3(in87, Not_Abus_3);
inv M2_Inv8_1_Inv4_0(in77, Not_Abus_4);
inv M2_Inv8_1_Inv4_1(in68, Not_Abus_5);
inv M2_Inv8_1_Inv4_2(in58, Not_Abus_6);
inv M2_Inv8_1_Inv4_3(in50, Not_Abus_7);
or2 M3_UM3_0_M8b3a_0_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_0_ContOr);
inv M3_UM3_0_M8b3a_0_Mux3a_1(in20, M3_UM3_0_M8b3a_0_NotContHi);
inv M3_UM3_0_M8b3a_0_Mux3a_2(M3_UM3_0_M8b3a_0_ContOr, M3_UM3_0_M8b3a_0_Cont00);
and2 M3_UM3_0_M8b3a_0_Mux3a_3(M3_UM3_0_M8b3a_0_NotContHi, M3_UM3_0_M8b3a_0_ContOr, M3_UM3_0_M8b3a_0_Cont01);
and2 M3_UM3_0_M8b3a_0_Mux3a_4(in97, M3_UM3_0_M8b3a_0_Cont00, M3_UM3_0_M8b3a_0_line4);
and2 M3_UM3_0_M8b3a_0_Mux3a_5(in283, M3_UM3_0_M8b3a_0_Cont01, M3_UM3_0_M8b3a_0_line5);
and2 M3_UM3_0_M8b3a_0_Mux3a_6(in116, in20, M3_UM3_0_M8b3a_0_line6);
or3 M3_UM3_0_M8b3a_0_Mux3a_7(M3_UM3_0_M8b3a_0_line4, M3_UM3_0_M8b3a_0_line5, M3_UM3_0_M8b3a_0_line6, M3_temp_0);
or2 M3_UM3_0_M8b3a_1_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_1_ContOr);
inv M3_UM3_0_M8b3a_1_Mux3a_1(in20, M3_UM3_0_M8b3a_1_NotContHi);
inv M3_UM3_0_M8b3a_1_Mux3a_2(M3_UM3_0_M8b3a_1_ContOr, M3_UM3_0_M8b3a_1_Cont00);
and2 M3_UM3_0_M8b3a_1_Mux3a_3(M3_UM3_0_M8b3a_1_NotContHi, M3_UM3_0_M8b3a_1_ContOr, M3_UM3_0_M8b3a_1_Cont01);
and2 M3_UM3_0_M8b3a_1_Mux3a_4(in87, M3_UM3_0_M8b3a_1_Cont00, M3_UM3_0_M8b3a_1_line4);
and2 M3_UM3_0_M8b3a_1_Mux3a_5(in116, M3_UM3_0_M8b3a_1_Cont01, M3_UM3_0_M8b3a_1_line5);
and2 M3_UM3_0_M8b3a_1_Mux3a_6(A_BCDbus_1, in20, M3_UM3_0_M8b3a_1_line6);
or3 M3_UM3_0_M8b3a_1_Mux3a_7(M3_UM3_0_M8b3a_1_line4, M3_UM3_0_M8b3a_1_line5, M3_UM3_0_M8b3a_1_line6, M3_temp_1);
or2 M3_UM3_0_M8b3a_2_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_2_ContOr);
inv M3_UM3_0_M8b3a_2_Mux3a_1(in20, M3_UM3_0_M8b3a_2_NotContHi);
inv M3_UM3_0_M8b3a_2_Mux3a_2(M3_UM3_0_M8b3a_2_ContOr, M3_UM3_0_M8b3a_2_Cont00);
and2 M3_UM3_0_M8b3a_2_Mux3a_3(M3_UM3_0_M8b3a_2_NotContHi, M3_UM3_0_M8b3a_2_ContOr, M3_UM3_0_M8b3a_2_Cont01);
and2 M3_UM3_0_M8b3a_2_Mux3a_4(in77, M3_UM3_0_M8b3a_2_Cont00, M3_UM3_0_M8b3a_2_line4);
and2 M3_UM3_0_M8b3a_2_Mux3a_5(in107, M3_UM3_0_M8b3a_2_Cont01, M3_UM3_0_M8b3a_2_line5);
and2 M3_UM3_0_M8b3a_2_Mux3a_6(A_BCDbus_2, in20, M3_UM3_0_M8b3a_2_line6);
or3 M3_UM3_0_M8b3a_2_Mux3a_7(M3_UM3_0_M8b3a_2_line4, M3_UM3_0_M8b3a_2_line5, M3_UM3_0_M8b3a_2_line6, M3_temp_2);
or2 M3_UM3_0_M8b3a_3_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_3_ContOr);
inv M3_UM3_0_M8b3a_3_Mux3a_1(in20, M3_UM3_0_M8b3a_3_NotContHi);
inv M3_UM3_0_M8b3a_3_Mux3a_2(M3_UM3_0_M8b3a_3_ContOr, M3_UM3_0_M8b3a_3_Cont00);
and2 M3_UM3_0_M8b3a_3_Mux3a_3(M3_UM3_0_M8b3a_3_NotContHi, M3_UM3_0_M8b3a_3_ContOr, M3_UM3_0_M8b3a_3_Cont01);
and2 M3_UM3_0_M8b3a_3_Mux3a_4(in68, M3_UM3_0_M8b3a_3_Cont00, M3_UM3_0_M8b3a_3_line4);
and2 M3_UM3_0_M8b3a_3_Mux3a_5(in97, M3_UM3_0_M8b3a_3_Cont01, M3_UM3_0_M8b3a_3_line5);
and2 M3_UM3_0_M8b3a_3_Mux3a_6(A_BCDbus_3, in20, M3_UM3_0_M8b3a_3_line6);
or3 M3_UM3_0_M8b3a_3_Mux3a_7(M3_UM3_0_M8b3a_3_line4, M3_UM3_0_M8b3a_3_line5, M3_UM3_0_M8b3a_3_line6, M3_temp_3);
or2 M3_UM3_0_M8b3a_4_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_4_ContOr);
inv M3_UM3_0_M8b3a_4_Mux3a_1(in20, M3_UM3_0_M8b3a_4_NotContHi);
inv M3_UM3_0_M8b3a_4_Mux3a_2(M3_UM3_0_M8b3a_4_ContOr, M3_UM3_0_M8b3a_4_Cont00);
and2 M3_UM3_0_M8b3a_4_Mux3a_3(M3_UM3_0_M8b3a_4_NotContHi, M3_UM3_0_M8b3a_4_ContOr, M3_UM3_0_M8b3a_4_Cont01);
and2 M3_UM3_0_M8b3a_4_Mux3a_4(in58, M3_UM3_0_M8b3a_4_Cont00, M3_UM3_0_M8b3a_4_line4);
and2 M3_UM3_0_M8b3a_4_Mux3a_5(in87, M3_UM3_0_M8b3a_4_Cont01, M3_UM3_0_M8b3a_4_line5);
and2 M3_UM3_0_M8b3a_4_Mux3a_6(in77, in20, M3_UM3_0_M8b3a_4_line6);
or3 M3_UM3_0_M8b3a_4_Mux3a_7(M3_UM3_0_M8b3a_4_line4, M3_UM3_0_M8b3a_4_line5, M3_UM3_0_M8b3a_4_line6, M3_temp_4);
or2 M3_UM3_0_M8b3a_5_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_5_ContOr);
inv M3_UM3_0_M8b3a_5_Mux3a_1(in20, M3_UM3_0_M8b3a_5_NotContHi);
inv M3_UM3_0_M8b3a_5_Mux3a_2(M3_UM3_0_M8b3a_5_ContOr, M3_UM3_0_M8b3a_5_Cont00);
and2 M3_UM3_0_M8b3a_5_Mux3a_3(M3_UM3_0_M8b3a_5_NotContHi, M3_UM3_0_M8b3a_5_ContOr, M3_UM3_0_M8b3a_5_Cont01);
and2 M3_UM3_0_M8b3a_5_Mux3a_4(in50, M3_UM3_0_M8b3a_5_Cont00, M3_UM3_0_M8b3a_5_line4);
and2 M3_UM3_0_M8b3a_5_Mux3a_5(in77, M3_UM3_0_M8b3a_5_Cont01, M3_UM3_0_M8b3a_5_line5);
and2 M3_UM3_0_M8b3a_5_Mux3a_6(A_BCDbus_5, in20, M3_UM3_0_M8b3a_5_line6);
or3 M3_UM3_0_M8b3a_5_Mux3a_7(M3_UM3_0_M8b3a_5_line4, M3_UM3_0_M8b3a_5_line5, M3_UM3_0_M8b3a_5_line6, M3_temp_5);
or2 M3_UM3_0_M8b3a_6_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_6_ContOr);
inv M3_UM3_0_M8b3a_6_Mux3a_1(in20, M3_UM3_0_M8b3a_6_NotContHi);
inv M3_UM3_0_M8b3a_6_Mux3a_2(M3_UM3_0_M8b3a_6_ContOr, M3_UM3_0_M8b3a_6_Cont00);
and2 M3_UM3_0_M8b3a_6_Mux3a_3(M3_UM3_0_M8b3a_6_NotContHi, M3_UM3_0_M8b3a_6_ContOr, M3_UM3_0_M8b3a_6_Cont01);
and2 M3_UM3_0_M8b3a_6_Mux3a_4(in159, M3_UM3_0_M8b3a_6_Cont00, M3_UM3_0_M8b3a_6_line4);
and2 M3_UM3_0_M8b3a_6_Mux3a_5(in68, M3_UM3_0_M8b3a_6_Cont01, M3_UM3_0_M8b3a_6_line5);
and2 M3_UM3_0_M8b3a_6_Mux3a_6(A_BCDbus_6, in20, M3_UM3_0_M8b3a_6_line6);
or3 M3_UM3_0_M8b3a_6_Mux3a_7(M3_UM3_0_M8b3a_6_line4, M3_UM3_0_M8b3a_6_line5, M3_UM3_0_M8b3a_6_line6, M3_temp_6);
or2 M3_UM3_0_M8b3a_7_Mux3a_0(in20, in33, M3_UM3_0_M8b3a_7_ContOr);
inv M3_UM3_0_M8b3a_7_Mux3a_1(in20, M3_UM3_0_M8b3a_7_NotContHi);
inv M3_UM3_0_M8b3a_7_Mux3a_2(M3_UM3_0_M8b3a_7_ContOr, M3_UM3_0_M8b3a_7_Cont00);
and2 M3_UM3_0_M8b3a_7_Mux3a_3(M3_UM3_0_M8b3a_7_NotContHi, M3_UM3_0_M8b3a_7_ContOr, M3_UM3_0_M8b3a_7_Cont01);
and2 M3_UM3_0_M8b3a_7_Mux3a_4(in150, M3_UM3_0_M8b3a_7_Cont00, M3_UM3_0_M8b3a_7_line4);
and2 M3_UM3_0_M8b3a_7_Mux3a_5(in58, M3_UM3_0_M8b3a_7_Cont01, M3_UM3_0_M8b3a_7_line5);
and2 M3_UM3_0_M8b3a_7_Mux3a_6(A_BCDbus_7, in20, M3_UM3_0_M8b3a_7_line6);
or3 M3_UM3_0_M8b3a_7_Mux3a_7(M3_UM3_0_M8b3a_7_line4, M3_UM3_0_M8b3a_7_line5, M3_UM3_0_M8b3a_7_line6, M3_temp_7);
nand2 M3_UM3_1(in1, in13, M3_line1);
nand3 M3_UM3_2(in1, in20, in33, M3_line2);
and2 M3_UM3_3(M3_line1, M3_line2, M3_line3);
inv M3_UM3_4(M3_line3, M3_MSel0);
and2 M3_UM3_5(in13, in20, M3_line5);
inv M3_UM3_6(M3_line5, M3_line6);
or2 M3_UM3_7(in1, M3_line6, M3_line7);
inv M3_UM3_8(M3_line7, M3_MSel2);
inv M3_UM3_9(in33, M3_line9);
inv M3_UM3_10(in20, M3_line10);
or2 M3_UM3_11(M3_line9, in1, M3_line11);
or2 M3_UM3_12(M3_line10, in1, M3_line12);
and3 M3_UM3_13(M3_line3, M3_line7, M3_line11, M3_MSel1a);
and3 M3_UM3_14(M3_line3, M3_line7, M3_line12, M3_MSel1b);
inv M3_UM3_15(M3_line11, M3_line15);
inv M3_UM3_16(M3_line12, M3_line16);
and3 M3_UM3_17(M3_line3, M3_line7, M3_line15, M3_MSel3a);
and3 M3_UM3_18(M3_line3, M3_line7, M3_line16, M3_MSel3b);
and2 M3_UM3_19_M4b4a_0_Mux4a_0(M3_temp_0, M3_MSel0, M3_UM3_19_M4b4a_0_line0);
and2 M3_UM3_19_M4b4a_0_Mux4a_1(in116, M3_MSel1a, M3_UM3_19_M4b4a_0_line1);
and2 M3_UM3_19_M4b4a_0_Mux4a_2(Not_Abus_0, M3_MSel2, M3_UM3_19_M4b4a_0_line2);
and2 M3_UM3_19_M4b4a_0_Mux4a_3(gnd, M3_MSel3a, M3_UM3_19_M4b4a_0_line3);
or4 M3_UM3_19_M4b4a_0_Mux4a_4(M3_UM3_19_M4b4a_0_line0, M3_UM3_19_M4b4a_0_line1, M3_UM3_19_M4b4a_0_line2, M3_UM3_19_M4b4a_0_line3, MAbus_0);
and2 M3_UM3_19_M4b4a_1_Mux4a_0(M3_temp_1, M3_MSel0, M3_UM3_19_M4b4a_1_line0);
and2 M3_UM3_19_M4b4a_1_Mux4a_1(in107, M3_MSel1a, M3_UM3_19_M4b4a_1_line1);
and2 M3_UM3_19_M4b4a_1_Mux4a_2(Not_Abus_1, M3_MSel2, M3_UM3_19_M4b4a_1_line2);
and2 M3_UM3_19_M4b4a_1_Mux4a_3(gnd, M3_MSel3a, M3_UM3_19_M4b4a_1_line3);
or4 M3_UM3_19_M4b4a_1_Mux4a_4(M3_UM3_19_M4b4a_1_line0, M3_UM3_19_M4b4a_1_line1, M3_UM3_19_M4b4a_1_line2, M3_UM3_19_M4b4a_1_line3, MAbus_1);
and2 M3_UM3_19_M4b4a_2_Mux4a_0(M3_temp_2, M3_MSel0, M3_UM3_19_M4b4a_2_line0);
and2 M3_UM3_19_M4b4a_2_Mux4a_1(in97, M3_MSel1a, M3_UM3_19_M4b4a_2_line1);
and2 M3_UM3_19_M4b4a_2_Mux4a_2(Not_Abus_2, M3_MSel2, M3_UM3_19_M4b4a_2_line2);
and2 M3_UM3_19_M4b4a_2_Mux4a_3(gnd, M3_MSel3a, M3_UM3_19_M4b4a_2_line3);
or4 M3_UM3_19_M4b4a_2_Mux4a_4(M3_UM3_19_M4b4a_2_line0, M3_UM3_19_M4b4a_2_line1, M3_UM3_19_M4b4a_2_line2, M3_UM3_19_M4b4a_2_line3, MAbus_2);
and2 M3_UM3_19_M4b4a_3_Mux4a_0(M3_temp_3, M3_MSel0, M3_UM3_19_M4b4a_3_line0);
and2 M3_UM3_19_M4b4a_3_Mux4a_1(in87, M3_MSel1a, M3_UM3_19_M4b4a_3_line1);
and2 M3_UM3_19_M4b4a_3_Mux4a_2(Not_Abus_3, M3_MSel2, M3_UM3_19_M4b4a_3_line2);
and2 M3_UM3_19_M4b4a_3_Mux4a_3(gnd, M3_MSel3a, M3_UM3_19_M4b4a_3_line3);
or4 M3_UM3_19_M4b4a_3_Mux4a_4(M3_UM3_19_M4b4a_3_line0, M3_UM3_19_M4b4a_3_line1, M3_UM3_19_M4b4a_3_line2, M3_UM3_19_M4b4a_3_line3, MAbus_3);
and2 M3_UM3_20_M4b4a_0_Mux4a_0(M3_temp_4, M3_MSel0, M3_UM3_20_M4b4a_0_line0);
and2 M3_UM3_20_M4b4a_0_Mux4a_1(in77, M3_MSel1b, M3_UM3_20_M4b4a_0_line1);
and2 M3_UM3_20_M4b4a_0_Mux4a_2(Not_Abus_4, M3_MSel2, M3_UM3_20_M4b4a_0_line2);
and2 M3_UM3_20_M4b4a_0_Mux4a_3(gnd, M3_MSel3b, M3_UM3_20_M4b4a_0_line3);
or4 M3_UM3_20_M4b4a_0_Mux4a_4(M3_UM3_20_M4b4a_0_line0, M3_UM3_20_M4b4a_0_line1, M3_UM3_20_M4b4a_0_line2, M3_UM3_20_M4b4a_0_line3, MAbus_4);
and2 M3_UM3_20_M4b4a_1_Mux4a_0(M3_temp_5, M3_MSel0, M3_UM3_20_M4b4a_1_line0);
and2 M3_UM3_20_M4b4a_1_Mux4a_1(in68, M3_MSel1b, M3_UM3_20_M4b4a_1_line1);
and2 M3_UM3_20_M4b4a_1_Mux4a_2(Not_Abus_5, M3_MSel2, M3_UM3_20_M4b4a_1_line2);
and2 M3_UM3_20_M4b4a_1_Mux4a_3(gnd, M3_MSel3b, M3_UM3_20_M4b4a_1_line3);
or4 M3_UM3_20_M4b4a_1_Mux4a_4(M3_UM3_20_M4b4a_1_line0, M3_UM3_20_M4b4a_1_line1, M3_UM3_20_M4b4a_1_line2, M3_UM3_20_M4b4a_1_line3, MAbus_5);
and2 M3_UM3_20_M4b4a_2_Mux4a_0(M3_temp_6, M3_MSel0, M3_UM3_20_M4b4a_2_line0);
and2 M3_UM3_20_M4b4a_2_Mux4a_1(in58, M3_MSel1b, M3_UM3_20_M4b4a_2_line1);
and2 M3_UM3_20_M4b4a_2_Mux4a_2(Not_Abus_6, M3_MSel2, M3_UM3_20_M4b4a_2_line2);
and2 M3_UM3_20_M4b4a_2_Mux4a_3(gnd, M3_MSel3b, M3_UM3_20_M4b4a_2_line3);
or4 M3_UM3_20_M4b4a_2_Mux4a_4(M3_UM3_20_M4b4a_2_line0, M3_UM3_20_M4b4a_2_line1, M3_UM3_20_M4b4a_2_line2, M3_UM3_20_M4b4a_2_line3, MAbus_6);
and2 M3_UM3_20_M4b4a_3_Mux4a_0(M3_temp_7, M3_MSel0, M3_UM3_20_M4b4a_3_line0);
and2 M3_UM3_20_M4b4a_3_Mux4a_1(in50, M3_MSel1b, M3_UM3_20_M4b4a_3_line1);
and2 M3_UM3_20_M4b4a_3_Mux4a_2(Not_Abus_7, M3_MSel2, M3_UM3_20_M4b4a_3_line2);
and2 M3_UM3_20_M4b4a_3_Mux4a_3(gnd, M3_MSel3b, M3_UM3_20_M4b4a_3_line3);
or4 M3_UM3_20_M4b4a_3_Mux4a_4(M3_UM3_20_M4b4a_3_line0, M3_UM3_20_M4b4a_3_line1, M3_UM3_20_M4b4a_3_line2, M3_UM3_20_M4b4a_3_line3, MAbus_7);
or2 M4_UM4_0_M8b3a_0_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_0_ContOr);
inv M4_UM4_0_M8b3a_0_Mux3a_1(in33, M4_UM4_0_M8b3a_0_NotContHi);
inv M4_UM4_0_M8b3a_0_Mux3a_2(M4_UM4_0_M8b3a_0_ContOr, M4_UM4_0_M8b3a_0_Cont00);
and2 M4_UM4_0_M8b3a_0_Mux3a_3(M4_UM4_0_M8b3a_0_NotContHi, M4_UM4_0_M8b3a_0_ContOr, M4_UM4_0_M8b3a_0_Cont01);
and2 M4_UM4_0_M8b3a_0_Mux3a_4(in257, M4_UM4_0_M8b3a_0_Cont00, M4_UM4_0_M8b3a_0_line4);
and2 M4_UM4_0_M8b3a_0_Mux3a_5(in264, M4_UM4_0_M8b3a_0_Cont01, M4_UM4_0_M8b3a_0_line5);
and2 M4_UM4_0_M8b3a_0_Mux3a_6(in303, in33, M4_UM4_0_M8b3a_0_line6);
or3 M4_UM4_0_M8b3a_0_Mux3a_7(M4_UM4_0_M8b3a_0_line4, M4_UM4_0_M8b3a_0_line5, M4_UM4_0_M8b3a_0_line6, M4_temp_0);
or2 M4_UM4_0_M8b3a_1_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_1_ContOr);
inv M4_UM4_0_M8b3a_1_Mux3a_1(in33, M4_UM4_0_M8b3a_1_NotContHi);
inv M4_UM4_0_M8b3a_1_Mux3a_2(M4_UM4_0_M8b3a_1_ContOr, M4_UM4_0_M8b3a_1_Cont00);
and2 M4_UM4_0_M8b3a_1_Mux3a_3(M4_UM4_0_M8b3a_1_NotContHi, M4_UM4_0_M8b3a_1_ContOr, M4_UM4_0_M8b3a_1_Cont01);
and2 M4_UM4_0_M8b3a_1_Mux3a_4(in250, M4_UM4_0_M8b3a_1_Cont00, M4_UM4_0_M8b3a_1_line4);
and2 M4_UM4_0_M8b3a_1_Mux3a_5(in257, M4_UM4_0_M8b3a_1_Cont01, M4_UM4_0_M8b3a_1_line5);
and2 M4_UM4_0_M8b3a_1_Mux3a_6(in294, in33, M4_UM4_0_M8b3a_1_line6);
or3 M4_UM4_0_M8b3a_1_Mux3a_7(M4_UM4_0_M8b3a_1_line4, M4_UM4_0_M8b3a_1_line5, M4_UM4_0_M8b3a_1_line6, M4_temp_1);
or2 M4_UM4_0_M8b3a_2_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_2_ContOr);
inv M4_UM4_0_M8b3a_2_Mux3a_1(in33, M4_UM4_0_M8b3a_2_NotContHi);
inv M4_UM4_0_M8b3a_2_Mux3a_2(M4_UM4_0_M8b3a_2_ContOr, M4_UM4_0_M8b3a_2_Cont00);
and2 M4_UM4_0_M8b3a_2_Mux3a_3(M4_UM4_0_M8b3a_2_NotContHi, M4_UM4_0_M8b3a_2_ContOr, M4_UM4_0_M8b3a_2_Cont01);
and2 M4_UM4_0_M8b3a_2_Mux3a_4(in244, M4_UM4_0_M8b3a_2_Cont00, M4_UM4_0_M8b3a_2_line4);
and2 M4_UM4_0_M8b3a_2_Mux3a_5(in250, M4_UM4_0_M8b3a_2_Cont01, M4_UM4_0_M8b3a_2_line5);
and2 M4_UM4_0_M8b3a_2_Mux3a_6(in283, in33, M4_UM4_0_M8b3a_2_line6);
or3 M4_UM4_0_M8b3a_2_Mux3a_7(M4_UM4_0_M8b3a_2_line4, M4_UM4_0_M8b3a_2_line5, M4_UM4_0_M8b3a_2_line6, M4_temp_2);
or2 M4_UM4_0_M8b3a_3_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_3_ContOr);
inv M4_UM4_0_M8b3a_3_Mux3a_1(in33, M4_UM4_0_M8b3a_3_NotContHi);
inv M4_UM4_0_M8b3a_3_Mux3a_2(M4_UM4_0_M8b3a_3_ContOr, M4_UM4_0_M8b3a_3_Cont00);
and2 M4_UM4_0_M8b3a_3_Mux3a_3(M4_UM4_0_M8b3a_3_NotContHi, M4_UM4_0_M8b3a_3_ContOr, M4_UM4_0_M8b3a_3_Cont01);
and2 M4_UM4_0_M8b3a_3_Mux3a_4(in238, M4_UM4_0_M8b3a_3_Cont00, M4_UM4_0_M8b3a_3_line4);
and2 M4_UM4_0_M8b3a_3_Mux3a_5(in244, M4_UM4_0_M8b3a_3_Cont01, M4_UM4_0_M8b3a_3_line5);
and2 M4_UM4_0_M8b3a_3_Mux3a_6(in116, in33, M4_UM4_0_M8b3a_3_line6);
or3 M4_UM4_0_M8b3a_3_Mux3a_7(M4_UM4_0_M8b3a_3_line4, M4_UM4_0_M8b3a_3_line5, M4_UM4_0_M8b3a_3_line6, M4_temp_3);
or2 M4_UM4_0_M8b3a_4_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_4_ContOr);
inv M4_UM4_0_M8b3a_4_Mux3a_1(in33, M4_UM4_0_M8b3a_4_NotContHi);
inv M4_UM4_0_M8b3a_4_Mux3a_2(M4_UM4_0_M8b3a_4_ContOr, M4_UM4_0_M8b3a_4_Cont00);
and2 M4_UM4_0_M8b3a_4_Mux3a_3(M4_UM4_0_M8b3a_4_NotContHi, M4_UM4_0_M8b3a_4_ContOr, M4_UM4_0_M8b3a_4_Cont01);
and2 M4_UM4_0_M8b3a_4_Mux3a_4(in232, M4_UM4_0_M8b3a_4_Cont00, M4_UM4_0_M8b3a_4_line4);
and2 M4_UM4_0_M8b3a_4_Mux3a_5(in238, M4_UM4_0_M8b3a_4_Cont01, M4_UM4_0_M8b3a_4_line5);
and2 M4_UM4_0_M8b3a_4_Mux3a_6(in107, in33, M4_UM4_0_M8b3a_4_line6);
or3 M4_UM4_0_M8b3a_4_Mux3a_7(M4_UM4_0_M8b3a_4_line4, M4_UM4_0_M8b3a_4_line5, M4_UM4_0_M8b3a_4_line6, M4_temp_4);
or2 M4_UM4_0_M8b3a_5_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_5_ContOr);
inv M4_UM4_0_M8b3a_5_Mux3a_1(in33, M4_UM4_0_M8b3a_5_NotContHi);
inv M4_UM4_0_M8b3a_5_Mux3a_2(M4_UM4_0_M8b3a_5_ContOr, M4_UM4_0_M8b3a_5_Cont00);
and2 M4_UM4_0_M8b3a_5_Mux3a_3(M4_UM4_0_M8b3a_5_NotContHi, M4_UM4_0_M8b3a_5_ContOr, M4_UM4_0_M8b3a_5_Cont01);
and2 M4_UM4_0_M8b3a_5_Mux3a_4(in226, M4_UM4_0_M8b3a_5_Cont00, M4_UM4_0_M8b3a_5_line4);
and2 M4_UM4_0_M8b3a_5_Mux3a_5(in232, M4_UM4_0_M8b3a_5_Cont01, M4_UM4_0_M8b3a_5_line5);
and2 M4_UM4_0_M8b3a_5_Mux3a_6(in97, in33, M4_UM4_0_M8b3a_5_line6);
or3 M4_UM4_0_M8b3a_5_Mux3a_7(M4_UM4_0_M8b3a_5_line4, M4_UM4_0_M8b3a_5_line5, M4_UM4_0_M8b3a_5_line6, M4_temp_5);
or2 M4_UM4_0_M8b3a_6_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_6_ContOr);
inv M4_UM4_0_M8b3a_6_Mux3a_1(in33, M4_UM4_0_M8b3a_6_NotContHi);
inv M4_UM4_0_M8b3a_6_Mux3a_2(M4_UM4_0_M8b3a_6_ContOr, M4_UM4_0_M8b3a_6_Cont00);
and2 M4_UM4_0_M8b3a_6_Mux3a_3(M4_UM4_0_M8b3a_6_NotContHi, M4_UM4_0_M8b3a_6_ContOr, M4_UM4_0_M8b3a_6_Cont01);
and2 M4_UM4_0_M8b3a_6_Mux3a_4(in223, M4_UM4_0_M8b3a_6_Cont00, M4_UM4_0_M8b3a_6_line4);
and2 M4_UM4_0_M8b3a_6_Mux3a_5(in226, M4_UM4_0_M8b3a_6_Cont01, M4_UM4_0_M8b3a_6_line5);
and2 M4_UM4_0_M8b3a_6_Mux3a_6(in87, in33, M4_UM4_0_M8b3a_6_line6);
or3 M4_UM4_0_M8b3a_6_Mux3a_7(M4_UM4_0_M8b3a_6_line4, M4_UM4_0_M8b3a_6_line5, M4_UM4_0_M8b3a_6_line6, M4_temp_6);
or2 M4_UM4_0_M8b3a_7_Mux3a_0(in33, in1698, M4_UM4_0_M8b3a_7_ContOr);
inv M4_UM4_0_M8b3a_7_Mux3a_1(in33, M4_UM4_0_M8b3a_7_NotContHi);
inv M4_UM4_0_M8b3a_7_Mux3a_2(M4_UM4_0_M8b3a_7_ContOr, M4_UM4_0_M8b3a_7_Cont00);
and2 M4_UM4_0_M8b3a_7_Mux3a_3(M4_UM4_0_M8b3a_7_NotContHi, M4_UM4_0_M8b3a_7_ContOr, M4_UM4_0_M8b3a_7_Cont01);
and2 M4_UM4_0_M8b3a_7_Mux3a_4(in222, M4_UM4_0_M8b3a_7_Cont00, M4_UM4_0_M8b3a_7_line4);
and2 M4_UM4_0_M8b3a_7_Mux3a_5(in223, M4_UM4_0_M8b3a_7_Cont01, M4_UM4_0_M8b3a_7_line5);
and2 M4_UM4_0_M8b3a_7_Mux3a_6(in77, in33, M4_UM4_0_M8b3a_7_line6);
or3 M4_UM4_0_M8b3a_7_Mux3a_7(M4_UM4_0_M8b3a_7_line4, M4_UM4_0_M8b3a_7_line5, M4_UM4_0_M8b3a_7_line6, M4_temp_7);
and2 M4_UM4_1(in33, in41, M4_line1);
inv M4_UM4_2(M4_line1, M4_line2);
and3 M4_UM4_3(in1, in13, M4_line2, M4_MSelHi);
inv M4_UM4_4(in1, M4_line4);
inv M4_UM4_5(in41, M4_line5);
and3 M4_UM4_6(M4_line4, in45, M4_line5, M4_MSelLo1);
and2 M4_UM4_7(M4_line4, in45, M4_MSelLo2);
or2 M4_UM4_8(in41, in45, M4_line8);
and2 M4_UM4_9(M4_line4, M4_line8, M4_MSelLo3);
inv M4_UM4_11_Mux3b_0(M4_MSelHi, M4_UM4_11_NotContHi);
inv M4_UM4_11_Mux3b_1(M4_MSelLo1, M4_UM4_11_NotContLo);
and3 M4_UM4_11_Mux3b_2(in270, M4_UM4_11_NotContHi, M4_UM4_11_NotContLo, M4_UM4_11_line2);
and3 M4_UM4_11_Mux3b_3(in274, M4_UM4_11_NotContHi, M4_MSelLo1, M4_UM4_11_line3);
and2 M4_UM4_11_Mux3b_4(M4_temp_0, M4_MSelHi, M4_UM4_11_line4);
or3 M4_UM4_11_Mux3b_5(M4_UM4_11_line2, M4_UM4_11_line3, M4_UM4_11_line4, MBbus_0);
inv M4_UM4_12_Mux3b_0(M4_MSelHi, M4_UM4_12_NotContHi);
inv M4_UM4_12_Mux3b_1(M4_MSelLo1, M4_UM4_12_NotContLo);
and3 M4_UM4_12_Mux3b_2(in264, M4_UM4_12_NotContHi, M4_UM4_12_NotContLo, M4_UM4_12_line2);
and3 M4_UM4_12_Mux3b_3(in274, M4_UM4_12_NotContHi, M4_MSelLo1, M4_UM4_12_line3);
and2 M4_UM4_12_Mux3b_4(M4_temp_1, M4_MSelHi, M4_UM4_12_line4);
or3 M4_UM4_12_Mux3b_5(M4_UM4_12_line2, M4_UM4_12_line3, M4_UM4_12_line4, MBbus_1);
inv M4_UM4_13_Mux3b_0(M4_MSelHi, M4_UM4_13_NotContHi);
inv M4_UM4_13_Mux3b_1(M4_MSelLo1, M4_UM4_13_NotContLo);
and3 M4_UM4_13_Mux3b_2(in257, M4_UM4_13_NotContHi, M4_UM4_13_NotContLo, M4_UM4_13_line2);
and3 M4_UM4_13_Mux3b_3(in274, M4_UM4_13_NotContHi, M4_MSelLo1, M4_UM4_13_line3);
and2 M4_UM4_13_Mux3b_4(M4_temp_2, M4_MSelHi, M4_UM4_13_line4);
or3 M4_UM4_13_Mux3b_5(M4_UM4_13_line2, M4_UM4_13_line3, M4_UM4_13_line4, MBbus_2);
inv M4_UM4_14_Mux3b_0(M4_MSelHi, M4_UM4_14_NotContHi);
inv M4_UM4_14_Mux3b_1(M4_MSelLo2, M4_UM4_14_NotContLo);
and3 M4_UM4_14_Mux3b_2(in250, M4_UM4_14_NotContHi, M4_UM4_14_NotContLo, M4_UM4_14_line2);
and3 M4_UM4_14_Mux3b_3(in274, M4_UM4_14_NotContHi, M4_MSelLo2, M4_UM4_14_line3);
and2 M4_UM4_14_Mux3b_4(M4_temp_3, M4_MSelHi, M4_UM4_14_line4);
or3 M4_UM4_14_Mux3b_5(M4_UM4_14_line2, M4_UM4_14_line3, M4_UM4_14_line4, MBbus_3);
inv M4_UM4_15_M4b3b_0_Mux3b_0(M4_MSelHi, M4_UM4_15_M4b3b_0_NotContHi);
inv M4_UM4_15_M4b3b_0_Mux3b_1(M4_MSelLo3, M4_UM4_15_M4b3b_0_NotContLo);
and3 M4_UM4_15_M4b3b_0_Mux3b_2(in244, M4_UM4_15_M4b3b_0_NotContHi, M4_UM4_15_M4b3b_0_NotContLo, M4_UM4_15_M4b3b_0_line2);
and3 M4_UM4_15_M4b3b_0_Mux3b_3(in274, M4_UM4_15_M4b3b_0_NotContHi, M4_MSelLo3, M4_UM4_15_M4b3b_0_line3);
and2 M4_UM4_15_M4b3b_0_Mux3b_4(M4_temp_4, M4_MSelHi, M4_UM4_15_M4b3b_0_line4);
or3 M4_UM4_15_M4b3b_0_Mux3b_5(M4_UM4_15_M4b3b_0_line2, M4_UM4_15_M4b3b_0_line3, M4_UM4_15_M4b3b_0_line4, MBbus_4);
inv M4_UM4_15_M4b3b_1_Mux3b_0(M4_MSelHi, M4_UM4_15_M4b3b_1_NotContHi);
inv M4_UM4_15_M4b3b_1_Mux3b_1(M4_MSelLo3, M4_UM4_15_M4b3b_1_NotContLo);
and3 M4_UM4_15_M4b3b_1_Mux3b_2(in238, M4_UM4_15_M4b3b_1_NotContHi, M4_UM4_15_M4b3b_1_NotContLo, M4_UM4_15_M4b3b_1_line2);
and3 M4_UM4_15_M4b3b_1_Mux3b_3(in274, M4_UM4_15_M4b3b_1_NotContHi, M4_MSelLo3, M4_UM4_15_M4b3b_1_line3);
and2 M4_UM4_15_M4b3b_1_Mux3b_4(M4_temp_5, M4_MSelHi, M4_UM4_15_M4b3b_1_line4);
or3 M4_UM4_15_M4b3b_1_Mux3b_5(M4_UM4_15_M4b3b_1_line2, M4_UM4_15_M4b3b_1_line3, M4_UM4_15_M4b3b_1_line4, MBbus_5);
inv M4_UM4_15_M4b3b_2_Mux3b_0(M4_MSelHi, M4_UM4_15_M4b3b_2_NotContHi);
inv M4_UM4_15_M4b3b_2_Mux3b_1(M4_MSelLo3, M4_UM4_15_M4b3b_2_NotContLo);
and3 M4_UM4_15_M4b3b_2_Mux3b_2(in232, M4_UM4_15_M4b3b_2_NotContHi, M4_UM4_15_M4b3b_2_NotContLo, M4_UM4_15_M4b3b_2_line2);
and3 M4_UM4_15_M4b3b_2_Mux3b_3(in274, M4_UM4_15_M4b3b_2_NotContHi, M4_MSelLo3, M4_UM4_15_M4b3b_2_line3);
and2 M4_UM4_15_M4b3b_2_Mux3b_4(M4_temp_6, M4_MSelHi, M4_UM4_15_M4b3b_2_line4);
or3 M4_UM4_15_M4b3b_2_Mux3b_5(M4_UM4_15_M4b3b_2_line2, M4_UM4_15_M4b3b_2_line3, M4_UM4_15_M4b3b_2_line4, MBbus_6);
inv M4_UM4_15_M4b3b_3_Mux3b_0(M4_MSelHi, M4_UM4_15_M4b3b_3_NotContHi);
inv M4_UM4_15_M4b3b_3_Mux3b_1(M4_MSelLo3, M4_UM4_15_M4b3b_3_NotContLo);
and3 M4_UM4_15_M4b3b_3_Mux3b_2(in226, M4_UM4_15_M4b3b_3_NotContHi, M4_UM4_15_M4b3b_3_NotContLo, M4_UM4_15_M4b3b_3_line2);
and3 M4_UM4_15_M4b3b_3_Mux3b_3(in274, M4_UM4_15_M4b3b_3_NotContHi, M4_MSelLo3, M4_UM4_15_M4b3b_3_line3);
and2 M4_UM4_15_M4b3b_3_Mux3b_4(M4_temp_7, M4_MSelHi, M4_UM4_15_M4b3b_3_line4);
or3 M4_UM4_15_M4b3b_3_Mux3b_5(M4_UM4_15_M4b3b_3_line2, M4_UM4_15_M4b3b_3_line3, M4_UM4_15_M4b3b_3_line4, MBbus_7);
inv M5_UM5_0(in1, M5_NotCont0);
inv M5_UM5_1(in20, M5_NotCont2);
and3 M5_UM5_2(M5_NotCont0, in13, M5_NotCont2, M5_ModeAux);
and3 M5_UM5_3(M5_ModeAux, in213, in343, M5_Mode);
and2 M5_UM5_4(M5_ModeAux, in213, M5_Mask7_6);
inv M5_UM5_5_LGP8_0_LGP0_Mux2_0(MBbus_0, M5_UM5_5_LGP8_0_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_0_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_0_LGP0_Not_ContIn, M5_UM5_5_LGP8_0_LGP0_line1);
and2 M5_UM5_5_LGP8_0_LGP0_Mux2_2(in200, MBbus_0, M5_UM5_5_LGP8_0_LGP0_line2);
or2 M5_UM5_5_LGP8_0_LGP0_Mux2_3(M5_UM5_5_LGP8_0_LGP0_line1, M5_UM5_5_LGP8_0_LGP0_line2, M5_UM5_5_LGP8_0_Mx0);
inv M5_UM5_5_LGP8_0_LGP1_Mux2_0(MBbus_0, M5_UM5_5_LGP8_0_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_0_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_0_LGP1_Not_ContIn, M5_UM5_5_LGP8_0_LGP1_line1);
and2 M5_UM5_5_LGP8_0_LGP1_Mux2_2(in169, MBbus_0, M5_UM5_5_LGP8_0_LGP1_line2);
or2 M5_UM5_5_LGP8_0_LGP1_Mux2_3(M5_UM5_5_LGP8_0_LGP1_line1, M5_UM5_5_LGP8_0_LGP1_line2, M5_UM5_5_LGP8_0_Mx1);
and2 M5_UM5_5_LGP8_0_LGP2(MAbus_0, M5_UM5_5_LGP8_0_Mx1, M5_Gbus_0);
or2 M5_UM5_5_LGP8_0_LGP3(MAbus_0, M5_UM5_5_LGP8_0_Mx0, M5_UM5_5_LGP8_0_InAMx0);
nand2 M5_UM5_5_LGP8_0_LGP4(MAbus_0, M5_UM5_5_LGP8_0_Mx1, M5_UM5_5_LGP8_0_InAMx1);
and2 M5_UM5_5_LGP8_0_LGP5(M5_UM5_5_LGP8_0_InAMx0, M5_UM5_5_LGP8_0_InAMx1, M5_Pbus_0);
and2 M5_UM5_5_LGP8_0_LGP6(M5_Mode, MAbus_0, M5_UM5_5_LGP8_0_InAMask);
inv M5_UM5_5_LGP8_0_LGP7_Xo0(M5_UM5_5_LGP8_0_InAMask, M5_UM5_5_LGP8_0_LGP7_NotA);
inv M5_UM5_5_LGP8_0_LGP7_Xo1(M5_Pbus_0, M5_UM5_5_LGP8_0_LGP7_NotB);
nand2 M5_UM5_5_LGP8_0_LGP7_Xo2(M5_UM5_5_LGP8_0_LGP7_NotA, M5_Pbus_0, M5_UM5_5_LGP8_0_LGP7_line2);
nand2 M5_UM5_5_LGP8_0_LGP7_Xo3(M5_UM5_5_LGP8_0_LGP7_NotB, M5_UM5_5_LGP8_0_InAMask, M5_UM5_5_LGP8_0_LGP7_line3);
nand2 M5_UM5_5_LGP8_0_LGP7_Xo4(M5_UM5_5_LGP8_0_LGP7_line2, M5_UM5_5_LGP8_0_LGP7_line3, XPbus_0);
inv M5_UM5_5_LGP8_0_LGP8(M5_Mode, M5_UM5_5_LGP8_0_NotMask);
and2 M5_UM5_5_LGP8_0_LGP9(M5_Gbus_0, M5_UM5_5_LGP8_0_NotMask, M5_XGbus_0);
inv M5_UM5_5_LGP8_1_LGP0_Mux2_0(MBbus_1, M5_UM5_5_LGP8_1_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_1_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_1_LGP0_Not_ContIn, M5_UM5_5_LGP8_1_LGP0_line1);
and2 M5_UM5_5_LGP8_1_LGP0_Mux2_2(in200, MBbus_1, M5_UM5_5_LGP8_1_LGP0_line2);
or2 M5_UM5_5_LGP8_1_LGP0_Mux2_3(M5_UM5_5_LGP8_1_LGP0_line1, M5_UM5_5_LGP8_1_LGP0_line2, M5_UM5_5_LGP8_1_Mx0);
inv M5_UM5_5_LGP8_1_LGP1_Mux2_0(MBbus_1, M5_UM5_5_LGP8_1_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_1_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_1_LGP1_Not_ContIn, M5_UM5_5_LGP8_1_LGP1_line1);
and2 M5_UM5_5_LGP8_1_LGP1_Mux2_2(in169, MBbus_1, M5_UM5_5_LGP8_1_LGP1_line2);
or2 M5_UM5_5_LGP8_1_LGP1_Mux2_3(M5_UM5_5_LGP8_1_LGP1_line1, M5_UM5_5_LGP8_1_LGP1_line2, M5_UM5_5_LGP8_1_Mx1);
and2 M5_UM5_5_LGP8_1_LGP2(MAbus_1, M5_UM5_5_LGP8_1_Mx1, M5_Gbus_1);
or2 M5_UM5_5_LGP8_1_LGP3(MAbus_1, M5_UM5_5_LGP8_1_Mx0, M5_UM5_5_LGP8_1_InAMx0);
nand2 M5_UM5_5_LGP8_1_LGP4(MAbus_1, M5_UM5_5_LGP8_1_Mx1, M5_UM5_5_LGP8_1_InAMx1);
and2 M5_UM5_5_LGP8_1_LGP5(M5_UM5_5_LGP8_1_InAMx0, M5_UM5_5_LGP8_1_InAMx1, M5_Pbus_1);
and2 M5_UM5_5_LGP8_1_LGP6(M5_Mode, MAbus_1, M5_UM5_5_LGP8_1_InAMask);
inv M5_UM5_5_LGP8_1_LGP7_Xo0(M5_UM5_5_LGP8_1_InAMask, M5_UM5_5_LGP8_1_LGP7_NotA);
inv M5_UM5_5_LGP8_1_LGP7_Xo1(M5_Pbus_1, M5_UM5_5_LGP8_1_LGP7_NotB);
nand2 M5_UM5_5_LGP8_1_LGP7_Xo2(M5_UM5_5_LGP8_1_LGP7_NotA, M5_Pbus_1, M5_UM5_5_LGP8_1_LGP7_line2);
nand2 M5_UM5_5_LGP8_1_LGP7_Xo3(M5_UM5_5_LGP8_1_LGP7_NotB, M5_UM5_5_LGP8_1_InAMask, M5_UM5_5_LGP8_1_LGP7_line3);
nand2 M5_UM5_5_LGP8_1_LGP7_Xo4(M5_UM5_5_LGP8_1_LGP7_line2, M5_UM5_5_LGP8_1_LGP7_line3, XPbus_1);
inv M5_UM5_5_LGP8_1_LGP8(M5_Mode, M5_UM5_5_LGP8_1_NotMask);
and2 M5_UM5_5_LGP8_1_LGP9(M5_Gbus_1, M5_UM5_5_LGP8_1_NotMask, M5_XGbus_1);
inv M5_UM5_5_LGP8_2_LGP0_Mux2_0(MBbus_2, M5_UM5_5_LGP8_2_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_2_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_2_LGP0_Not_ContIn, M5_UM5_5_LGP8_2_LGP0_line1);
and2 M5_UM5_5_LGP8_2_LGP0_Mux2_2(in200, MBbus_2, M5_UM5_5_LGP8_2_LGP0_line2);
or2 M5_UM5_5_LGP8_2_LGP0_Mux2_3(M5_UM5_5_LGP8_2_LGP0_line1, M5_UM5_5_LGP8_2_LGP0_line2, M5_UM5_5_LGP8_2_Mx0);
inv M5_UM5_5_LGP8_2_LGP1_Mux2_0(MBbus_2, M5_UM5_5_LGP8_2_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_2_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_2_LGP1_Not_ContIn, M5_UM5_5_LGP8_2_LGP1_line1);
and2 M5_UM5_5_LGP8_2_LGP1_Mux2_2(in169, MBbus_2, M5_UM5_5_LGP8_2_LGP1_line2);
or2 M5_UM5_5_LGP8_2_LGP1_Mux2_3(M5_UM5_5_LGP8_2_LGP1_line1, M5_UM5_5_LGP8_2_LGP1_line2, M5_UM5_5_LGP8_2_Mx1);
and2 M5_UM5_5_LGP8_2_LGP2(MAbus_2, M5_UM5_5_LGP8_2_Mx1, M5_Gbus_2);
or2 M5_UM5_5_LGP8_2_LGP3(MAbus_2, M5_UM5_5_LGP8_2_Mx0, M5_UM5_5_LGP8_2_InAMx0);
nand2 M5_UM5_5_LGP8_2_LGP4(MAbus_2, M5_UM5_5_LGP8_2_Mx1, M5_UM5_5_LGP8_2_InAMx1);
and2 M5_UM5_5_LGP8_2_LGP5(M5_UM5_5_LGP8_2_InAMx0, M5_UM5_5_LGP8_2_InAMx1, M5_Pbus_2);
and2 M5_UM5_5_LGP8_2_LGP6(M5_Mode, MAbus_2, M5_UM5_5_LGP8_2_InAMask);
inv M5_UM5_5_LGP8_2_LGP7_Xo0(M5_UM5_5_LGP8_2_InAMask, M5_UM5_5_LGP8_2_LGP7_NotA);
inv M5_UM5_5_LGP8_2_LGP7_Xo1(M5_Pbus_2, M5_UM5_5_LGP8_2_LGP7_NotB);
nand2 M5_UM5_5_LGP8_2_LGP7_Xo2(M5_UM5_5_LGP8_2_LGP7_NotA, M5_Pbus_2, M5_UM5_5_LGP8_2_LGP7_line2);
nand2 M5_UM5_5_LGP8_2_LGP7_Xo3(M5_UM5_5_LGP8_2_LGP7_NotB, M5_UM5_5_LGP8_2_InAMask, M5_UM5_5_LGP8_2_LGP7_line3);
nand2 M5_UM5_5_LGP8_2_LGP7_Xo4(M5_UM5_5_LGP8_2_LGP7_line2, M5_UM5_5_LGP8_2_LGP7_line3, XPbus_2);
inv M5_UM5_5_LGP8_2_LGP8(M5_Mode, M5_UM5_5_LGP8_2_NotMask);
and2 M5_UM5_5_LGP8_2_LGP9(M5_Gbus_2, M5_UM5_5_LGP8_2_NotMask, M5_XGbus_2);
inv M5_UM5_5_LGP8_3_LGP0_Mux2_0(MBbus_3, M5_UM5_5_LGP8_3_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_3_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_3_LGP0_Not_ContIn, M5_UM5_5_LGP8_3_LGP0_line1);
and2 M5_UM5_5_LGP8_3_LGP0_Mux2_2(in200, MBbus_3, M5_UM5_5_LGP8_3_LGP0_line2);
or2 M5_UM5_5_LGP8_3_LGP0_Mux2_3(M5_UM5_5_LGP8_3_LGP0_line1, M5_UM5_5_LGP8_3_LGP0_line2, M5_UM5_5_LGP8_3_Mx0);
inv M5_UM5_5_LGP8_3_LGP1_Mux2_0(MBbus_3, M5_UM5_5_LGP8_3_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_3_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_3_LGP1_Not_ContIn, M5_UM5_5_LGP8_3_LGP1_line1);
and2 M5_UM5_5_LGP8_3_LGP1_Mux2_2(in169, MBbus_3, M5_UM5_5_LGP8_3_LGP1_line2);
or2 M5_UM5_5_LGP8_3_LGP1_Mux2_3(M5_UM5_5_LGP8_3_LGP1_line1, M5_UM5_5_LGP8_3_LGP1_line2, M5_UM5_5_LGP8_3_Mx1);
and2 M5_UM5_5_LGP8_3_LGP2(MAbus_3, M5_UM5_5_LGP8_3_Mx1, M5_Gbus_3);
or2 M5_UM5_5_LGP8_3_LGP3(MAbus_3, M5_UM5_5_LGP8_3_Mx0, M5_UM5_5_LGP8_3_InAMx0);
nand2 M5_UM5_5_LGP8_3_LGP4(MAbus_3, M5_UM5_5_LGP8_3_Mx1, M5_UM5_5_LGP8_3_InAMx1);
and2 M5_UM5_5_LGP8_3_LGP5(M5_UM5_5_LGP8_3_InAMx0, M5_UM5_5_LGP8_3_InAMx1, M5_Pbus_3);
and2 M5_UM5_5_LGP8_3_LGP6(M5_Mode, MAbus_3, M5_UM5_5_LGP8_3_InAMask);
inv M5_UM5_5_LGP8_3_LGP7_Xo0(M5_UM5_5_LGP8_3_InAMask, M5_UM5_5_LGP8_3_LGP7_NotA);
inv M5_UM5_5_LGP8_3_LGP7_Xo1(M5_Pbus_3, M5_UM5_5_LGP8_3_LGP7_NotB);
nand2 M5_UM5_5_LGP8_3_LGP7_Xo2(M5_UM5_5_LGP8_3_LGP7_NotA, M5_Pbus_3, M5_UM5_5_LGP8_3_LGP7_line2);
nand2 M5_UM5_5_LGP8_3_LGP7_Xo3(M5_UM5_5_LGP8_3_LGP7_NotB, M5_UM5_5_LGP8_3_InAMask, M5_UM5_5_LGP8_3_LGP7_line3);
nand2 M5_UM5_5_LGP8_3_LGP7_Xo4(M5_UM5_5_LGP8_3_LGP7_line2, M5_UM5_5_LGP8_3_LGP7_line3, XPbus_3);
inv M5_UM5_5_LGP8_3_LGP8(M5_Mode, M5_UM5_5_LGP8_3_NotMask);
and2 M5_UM5_5_LGP8_3_LGP9(M5_Gbus_3, M5_UM5_5_LGP8_3_NotMask, M5_XGbus_3);
inv M5_UM5_5_LGP8_4_LGP0_Mux2_0(MBbus_4, M5_UM5_5_LGP8_4_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_4_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_4_LGP0_Not_ContIn, M5_UM5_5_LGP8_4_LGP0_line1);
and2 M5_UM5_5_LGP8_4_LGP0_Mux2_2(in200, MBbus_4, M5_UM5_5_LGP8_4_LGP0_line2);
or2 M5_UM5_5_LGP8_4_LGP0_Mux2_3(M5_UM5_5_LGP8_4_LGP0_line1, M5_UM5_5_LGP8_4_LGP0_line2, M5_UM5_5_LGP8_4_Mx0);
inv M5_UM5_5_LGP8_4_LGP1_Mux2_0(MBbus_4, M5_UM5_5_LGP8_4_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_4_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_4_LGP1_Not_ContIn, M5_UM5_5_LGP8_4_LGP1_line1);
and2 M5_UM5_5_LGP8_4_LGP1_Mux2_2(in169, MBbus_4, M5_UM5_5_LGP8_4_LGP1_line2);
or2 M5_UM5_5_LGP8_4_LGP1_Mux2_3(M5_UM5_5_LGP8_4_LGP1_line1, M5_UM5_5_LGP8_4_LGP1_line2, M5_UM5_5_LGP8_4_Mx1);
and2 M5_UM5_5_LGP8_4_LGP2(MAbus_4, M5_UM5_5_LGP8_4_Mx1, M5_Gbus_4);
or2 M5_UM5_5_LGP8_4_LGP3(MAbus_4, M5_UM5_5_LGP8_4_Mx0, M5_UM5_5_LGP8_4_InAMx0);
nand2 M5_UM5_5_LGP8_4_LGP4(MAbus_4, M5_UM5_5_LGP8_4_Mx1, M5_UM5_5_LGP8_4_InAMx1);
and2 M5_UM5_5_LGP8_4_LGP5(M5_UM5_5_LGP8_4_InAMx0, M5_UM5_5_LGP8_4_InAMx1, M5_Pbus_4);
and2 M5_UM5_5_LGP8_4_LGP6(M5_Mode, MAbus_4, M5_UM5_5_LGP8_4_InAMask);
inv M5_UM5_5_LGP8_4_LGP7_Xo0(M5_UM5_5_LGP8_4_InAMask, M5_UM5_5_LGP8_4_LGP7_NotA);
inv M5_UM5_5_LGP8_4_LGP7_Xo1(M5_Pbus_4, M5_UM5_5_LGP8_4_LGP7_NotB);
nand2 M5_UM5_5_LGP8_4_LGP7_Xo2(M5_UM5_5_LGP8_4_LGP7_NotA, M5_Pbus_4, M5_UM5_5_LGP8_4_LGP7_line2);
nand2 M5_UM5_5_LGP8_4_LGP7_Xo3(M5_UM5_5_LGP8_4_LGP7_NotB, M5_UM5_5_LGP8_4_InAMask, M5_UM5_5_LGP8_4_LGP7_line3);
nand2 M5_UM5_5_LGP8_4_LGP7_Xo4(M5_UM5_5_LGP8_4_LGP7_line2, M5_UM5_5_LGP8_4_LGP7_line3, XPbus_4);
inv M5_UM5_5_LGP8_4_LGP8(M5_Mode, M5_UM5_5_LGP8_4_NotMask);
and2 M5_UM5_5_LGP8_4_LGP9(M5_Gbus_4, M5_UM5_5_LGP8_4_NotMask, M5_XGbus_4);
inv M5_UM5_5_LGP8_5_LGP0_Mux2_0(MBbus_5, M5_UM5_5_LGP8_5_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_5_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_5_LGP0_Not_ContIn, M5_UM5_5_LGP8_5_LGP0_line1);
and2 M5_UM5_5_LGP8_5_LGP0_Mux2_2(in200, MBbus_5, M5_UM5_5_LGP8_5_LGP0_line2);
or2 M5_UM5_5_LGP8_5_LGP0_Mux2_3(M5_UM5_5_LGP8_5_LGP0_line1, M5_UM5_5_LGP8_5_LGP0_line2, M5_UM5_5_LGP8_5_Mx0);
inv M5_UM5_5_LGP8_5_LGP1_Mux2_0(MBbus_5, M5_UM5_5_LGP8_5_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_5_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_5_LGP1_Not_ContIn, M5_UM5_5_LGP8_5_LGP1_line1);
and2 M5_UM5_5_LGP8_5_LGP1_Mux2_2(in169, MBbus_5, M5_UM5_5_LGP8_5_LGP1_line2);
or2 M5_UM5_5_LGP8_5_LGP1_Mux2_3(M5_UM5_5_LGP8_5_LGP1_line1, M5_UM5_5_LGP8_5_LGP1_line2, M5_UM5_5_LGP8_5_Mx1);
and2 M5_UM5_5_LGP8_5_LGP2(MAbus_5, M5_UM5_5_LGP8_5_Mx1, M5_Gbus_5);
or2 M5_UM5_5_LGP8_5_LGP3(MAbus_5, M5_UM5_5_LGP8_5_Mx0, M5_UM5_5_LGP8_5_InAMx0);
nand2 M5_UM5_5_LGP8_5_LGP4(MAbus_5, M5_UM5_5_LGP8_5_Mx1, M5_UM5_5_LGP8_5_InAMx1);
and2 M5_UM5_5_LGP8_5_LGP5(M5_UM5_5_LGP8_5_InAMx0, M5_UM5_5_LGP8_5_InAMx1, M5_Pbus_5);
and2 M5_UM5_5_LGP8_5_LGP6(M5_Mode, MAbus_5, M5_UM5_5_LGP8_5_InAMask);
inv M5_UM5_5_LGP8_5_LGP7_Xo0(M5_UM5_5_LGP8_5_InAMask, M5_UM5_5_LGP8_5_LGP7_NotA);
inv M5_UM5_5_LGP8_5_LGP7_Xo1(M5_Pbus_5, M5_UM5_5_LGP8_5_LGP7_NotB);
nand2 M5_UM5_5_LGP8_5_LGP7_Xo2(M5_UM5_5_LGP8_5_LGP7_NotA, M5_Pbus_5, M5_UM5_5_LGP8_5_LGP7_line2);
nand2 M5_UM5_5_LGP8_5_LGP7_Xo3(M5_UM5_5_LGP8_5_LGP7_NotB, M5_UM5_5_LGP8_5_InAMask, M5_UM5_5_LGP8_5_LGP7_line3);
nand2 M5_UM5_5_LGP8_5_LGP7_Xo4(M5_UM5_5_LGP8_5_LGP7_line2, M5_UM5_5_LGP8_5_LGP7_line3, XPbus_5);
inv M5_UM5_5_LGP8_5_LGP8(M5_Mode, M5_UM5_5_LGP8_5_NotMask);
and2 M5_UM5_5_LGP8_5_LGP9(M5_Gbus_5, M5_UM5_5_LGP8_5_NotMask, M5_XGbus_5);
inv M5_UM5_5_LGP8_6_LGP0_Mux2_0(MBbus_6, M5_UM5_5_LGP8_6_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_6_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_6_LGP0_Not_ContIn, M5_UM5_5_LGP8_6_LGP0_line1);
and2 M5_UM5_5_LGP8_6_LGP0_Mux2_2(in200, MBbus_6, M5_UM5_5_LGP8_6_LGP0_line2);
or2 M5_UM5_5_LGP8_6_LGP0_Mux2_3(M5_UM5_5_LGP8_6_LGP0_line1, M5_UM5_5_LGP8_6_LGP0_line2, M5_UM5_5_LGP8_6_Mx0);
inv M5_UM5_5_LGP8_6_LGP1_Mux2_0(MBbus_6, M5_UM5_5_LGP8_6_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_6_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_6_LGP1_Not_ContIn, M5_UM5_5_LGP8_6_LGP1_line1);
and2 M5_UM5_5_LGP8_6_LGP1_Mux2_2(in169, MBbus_6, M5_UM5_5_LGP8_6_LGP1_line2);
or2 M5_UM5_5_LGP8_6_LGP1_Mux2_3(M5_UM5_5_LGP8_6_LGP1_line1, M5_UM5_5_LGP8_6_LGP1_line2, M5_UM5_5_LGP8_6_Mx1);
and2 M5_UM5_5_LGP8_6_LGP2(MAbus_6, M5_UM5_5_LGP8_6_Mx1, M5_Gbus_6);
or2 M5_UM5_5_LGP8_6_LGP3(MAbus_6, M5_UM5_5_LGP8_6_Mx0, M5_UM5_5_LGP8_6_InAMx0);
nand2 M5_UM5_5_LGP8_6_LGP4(MAbus_6, M5_UM5_5_LGP8_6_Mx1, M5_UM5_5_LGP8_6_InAMx1);
and2 M5_UM5_5_LGP8_6_LGP5(M5_UM5_5_LGP8_6_InAMx0, M5_UM5_5_LGP8_6_InAMx1, M5_Pbus_6);
and2 M5_UM5_5_LGP8_6_LGP6(M5_Mask7_6, MAbus_6, M5_UM5_5_LGP8_6_InAMask);
inv M5_UM5_5_LGP8_6_LGP7_Xo0(M5_UM5_5_LGP8_6_InAMask, M5_UM5_5_LGP8_6_LGP7_NotA);
inv M5_UM5_5_LGP8_6_LGP7_Xo1(M5_Pbus_6, M5_UM5_5_LGP8_6_LGP7_NotB);
nand2 M5_UM5_5_LGP8_6_LGP7_Xo2(M5_UM5_5_LGP8_6_LGP7_NotA, M5_Pbus_6, M5_UM5_5_LGP8_6_LGP7_line2);
nand2 M5_UM5_5_LGP8_6_LGP7_Xo3(M5_UM5_5_LGP8_6_LGP7_NotB, M5_UM5_5_LGP8_6_InAMask, M5_UM5_5_LGP8_6_LGP7_line3);
nand2 M5_UM5_5_LGP8_6_LGP7_Xo4(M5_UM5_5_LGP8_6_LGP7_line2, M5_UM5_5_LGP8_6_LGP7_line3, XPbus_6);
inv M5_UM5_5_LGP8_6_LGP8(M5_Mask7_6, M5_UM5_5_LGP8_6_NotMask);
and2 M5_UM5_5_LGP8_6_LGP9(M5_Gbus_6, M5_UM5_5_LGP8_6_NotMask, M5_XGbus_6);
inv M5_UM5_5_LGP8_7_LGP0_Mux2_0(MBbus_7, M5_UM5_5_LGP8_7_LGP0_Not_ContIn);
and2 M5_UM5_5_LGP8_7_LGP0_Mux2_1(in190, M5_UM5_5_LGP8_7_LGP0_Not_ContIn, M5_UM5_5_LGP8_7_LGP0_line1);
and2 M5_UM5_5_LGP8_7_LGP0_Mux2_2(in200, MBbus_7, M5_UM5_5_LGP8_7_LGP0_line2);
or2 M5_UM5_5_LGP8_7_LGP0_Mux2_3(M5_UM5_5_LGP8_7_LGP0_line1, M5_UM5_5_LGP8_7_LGP0_line2, M5_UM5_5_LGP8_7_Mx0);
inv M5_UM5_5_LGP8_7_LGP1_Mux2_0(MBbus_7, M5_UM5_5_LGP8_7_LGP1_Not_ContIn);
and2 M5_UM5_5_LGP8_7_LGP1_Mux2_1(in179, M5_UM5_5_LGP8_7_LGP1_Not_ContIn, M5_UM5_5_LGP8_7_LGP1_line1);
and2 M5_UM5_5_LGP8_7_LGP1_Mux2_2(in169, MBbus_7, M5_UM5_5_LGP8_7_LGP1_line2);
or2 M5_UM5_5_LGP8_7_LGP1_Mux2_3(M5_UM5_5_LGP8_7_LGP1_line1, M5_UM5_5_LGP8_7_LGP1_line2, M5_UM5_5_LGP8_7_Mx1);
and2 M5_UM5_5_LGP8_7_LGP2(MAbus_7, M5_UM5_5_LGP8_7_Mx1, M5_Gbus_7);
or2 M5_UM5_5_LGP8_7_LGP3(MAbus_7, M5_UM5_5_LGP8_7_Mx0, M5_UM5_5_LGP8_7_InAMx0);
nand2 M5_UM5_5_LGP8_7_LGP4(MAbus_7, M5_UM5_5_LGP8_7_Mx1, M5_UM5_5_LGP8_7_InAMx1);
and2 M5_UM5_5_LGP8_7_LGP5(M5_UM5_5_LGP8_7_InAMx0, M5_UM5_5_LGP8_7_InAMx1, M5_Pbus_7);
and2 M5_UM5_5_LGP8_7_LGP6(M5_Mask7_6, MAbus_7, M5_UM5_5_LGP8_7_InAMask);
inv M5_UM5_5_LGP8_7_LGP7_Xo0(M5_UM5_5_LGP8_7_InAMask, M5_UM5_5_LGP8_7_LGP7_NotA);
inv M5_UM5_5_LGP8_7_LGP7_Xo1(M5_Pbus_7, M5_UM5_5_LGP8_7_LGP7_NotB);
nand2 M5_UM5_5_LGP8_7_LGP7_Xo2(M5_UM5_5_LGP8_7_LGP7_NotA, M5_Pbus_7, M5_UM5_5_LGP8_7_LGP7_line2);
nand2 M5_UM5_5_LGP8_7_LGP7_Xo3(M5_UM5_5_LGP8_7_LGP7_NotB, M5_UM5_5_LGP8_7_InAMask, M5_UM5_5_LGP8_7_LGP7_line3);
nand2 M5_UM5_5_LGP8_7_LGP7_Xo4(M5_UM5_5_LGP8_7_LGP7_line2, M5_UM5_5_LGP8_7_LGP7_line3, XPbus_7);
inv M5_UM5_5_LGP8_7_LGP8(M5_Mask7_6, M5_UM5_5_LGP8_7_NotMask);
and2 M5_UM5_5_LGP8_7_LGP9(M5_Gbus_7, M5_UM5_5_LGP8_7_NotMask, M5_XGbus_7);
and4 M5_UM5_6_CC0(M5_Pbus_0, M5_Pbus_1, M5_Pbus_2, M5_Pbus_3, M5_UM5_6_PropLo);
and4 M5_UM5_6_CC1(M5_Pbus_4, M5_Pbus_5, M5_Pbus_6, M5_Pbus_7, M5_UM5_6_PropHi);
and2 M5_UM5_6_CC2(M5_UM5_6_PropLo, M5_UM5_6_PropHi, out372);
inv M5_UM5_6_CC3(M5_Mode, M5_UM5_6_NotMode);
and4 M5_UM5_6_CC4_CCP0(MBbus_0, MBbus_1, MBbus_2, MBbus_3, M5_UM5_6_CC4_InBLoAND);
nor4 M5_UM5_6_CC4_CCP1(MBbus_0, MBbus_1, MBbus_2, MBbus_3, M5_UM5_6_CC4_InBLoNOR);
inv M5_UM5_6_CC4_CCP2_Mux2_0(in179, M5_UM5_6_CC4_CCP2_Not_ContIn);
and2 M5_UM5_6_CC4_CCP2_Mux2_1(M5_UM5_6_CC4_InBLoAND, M5_UM5_6_CC4_CCP2_Not_ContIn, M5_UM5_6_CC4_CCP2_line1);
and2 M5_UM5_6_CC4_CCP2_Mux2_2(M5_UM5_6_CC4_InBLoNOR, in179, M5_UM5_6_CC4_CCP2_line2);
or2 M5_UM5_6_CC4_CCP2_Mux2_3(M5_UM5_6_CC4_CCP2_line1, M5_UM5_6_CC4_CCP2_line2, M5_UM5_6_CC4_InBprop);
inv M5_UM5_6_CC4_CCP3_Mux2_0(M5_Mode, M5_UM5_6_CC4_CCP3_Not_ContIn);
and2 M5_UM5_6_CC4_CCP3_Mux2_1(M5_UM5_6_PropLo, M5_UM5_6_CC4_CCP3_Not_ContIn, M5_UM5_6_CC4_CCP3_line1);
and2 M5_UM5_6_CC4_CCP3_Mux2_2(M5_UM5_6_CC4_InBprop, M5_Mode, M5_UM5_6_CC4_CCP3_line2);
or2 M5_UM5_6_CC4_CCP3_Mux2_3(M5_UM5_6_CC4_CCP3_line1, M5_UM5_6_CC4_CCP3_line2, M5_UM5_6_CC4_Pr);
and2 M5_UM5_6_CC4_CCP4(in330, M5_UM5_6_CC4_Pr, M5_UM5_6_CinPropLo);
and2 M5_UM5_6_CC5_Ao4a_0(M5_Pbus_3, M5_Gbus_2, M5_UM5_6_CC5_line0);
and3 M5_UM5_6_CC5_Ao4a_1(M5_Pbus_3, M5_Pbus_2, M5_Gbus_1, M5_UM5_6_CC5_line1);
and4 M5_UM5_6_CC5_Ao4a_2(M5_Pbus_3, M5_Pbus_2, M5_Pbus_1, M5_Gbus_0, M5_UM5_6_CC5_line2);
or4 M5_UM5_6_CC5_Ao4a_3(M5_Gbus_3, M5_UM5_6_CC5_line0, M5_UM5_6_CC5_line1, M5_UM5_6_CC5_line2, M5_UM5_6_LocalC0Lo);
and2 M5_UM5_6_CC6_Ao4a_0(M5_Pbus_7, M5_Gbus_6, M5_UM5_6_CC6_line0);
and3 M5_UM5_6_CC6_Ao4a_1(M5_Pbus_7, M5_Pbus_6, M5_Gbus_5, M5_UM5_6_CC6_line1);
and4 M5_UM5_6_CC6_Ao4a_2(M5_Pbus_7, M5_Pbus_6, M5_Pbus_5, M5_Gbus_4, M5_UM5_6_CC6_line2);
or4 M5_UM5_6_CC6_Ao4a_3(M5_Gbus_7, M5_UM5_6_CC6_line0, M5_UM5_6_CC6_line1, M5_UM5_6_CC6_line2, M5_UM5_6_LocalC0Hi);
and2 M5_UM5_6_CC7(M5_UM5_6_LocalC0Lo, M5_UM5_6_NotMode, M5_UM5_6_LoC0_M);
and2 M5_UM5_6_CC8_Cb0_Cla4_0_Ao2_0(XPbus_0, gnd, M5_UM5_6_CC8_Cb0_Cla4_0_line0);
or2 M5_UM5_6_CC8_Cb0_Cla4_0_Ao2_1(M5_XGbus_0, M5_UM5_6_CC8_Cb0_Cla4_0_line0, M5_UM5_6_CC8_Cy1bus_1);
and2 M5_UM5_6_CC8_Cb0_Cla4_1_Ao3a_0(XPbus_1, M5_XGbus_0, M5_UM5_6_CC8_Cb0_Cla4_1_line0);
and3 M5_UM5_6_CC8_Cb0_Cla4_1_Ao3a_1(XPbus_1, XPbus_0, gnd, M5_UM5_6_CC8_Cb0_Cla4_1_line1);
or3 M5_UM5_6_CC8_Cb0_Cla4_1_Ao3a_2(M5_XGbus_1, M5_UM5_6_CC8_Cb0_Cla4_1_line0, M5_UM5_6_CC8_Cb0_Cla4_1_line1, M5_UM5_6_CC8_Cy1bus_2);
and2 M5_UM5_6_CC8_Cb0_Cla4_2_Ao4a_0(XPbus_2, M5_XGbus_1, M5_UM5_6_CC8_Cb0_Cla4_2_line0);
and3 M5_UM5_6_CC8_Cb0_Cla4_2_Ao4a_1(XPbus_2, XPbus_1, M5_XGbus_0, M5_UM5_6_CC8_Cb0_Cla4_2_line1);
and4 M5_UM5_6_CC8_Cb0_Cla4_2_Ao4a_2(XPbus_2, XPbus_1, XPbus_0, gnd, M5_UM5_6_CC8_Cb0_Cla4_2_line2);
or4 M5_UM5_6_CC8_Cb0_Cla4_2_Ao4a_3(M5_XGbus_2, M5_UM5_6_CC8_Cb0_Cla4_2_line0, M5_UM5_6_CC8_Cb0_Cla4_2_line1, M5_UM5_6_CC8_Cb0_Cla4_2_line2, M5_UM5_6_CC8_Cy1bus_3);
and2 M5_UM5_6_CC8_Cb1_CP0(XPbus_0, in330, M5_UM5_6_CC8_Cy2bus_1);
and3 M5_UM5_6_CC8_Cb1_CP1(XPbus_1, XPbus_0, in330, M5_UM5_6_CC8_Cy2bus_2);
and4 M5_UM5_6_CC8_Cb1_CP2(XPbus_2, XPbus_1, XPbus_0, in330, M5_UM5_6_CC8_Cy2bus_3);
inv M5_UM5_6_CC8_Cb2_X4_0_Xo0(gnd, M5_UM5_6_CC8_Cb2_X4_0_NotA);
inv M5_UM5_6_CC8_Cb2_X4_0_Xo1(in330, M5_UM5_6_CC8_Cb2_X4_0_NotB);
nand2 M5_UM5_6_CC8_Cb2_X4_0_Xo2(M5_UM5_6_CC8_Cb2_X4_0_NotA, in330, M5_UM5_6_CC8_Cb2_X4_0_line2);
nand2 M5_UM5_6_CC8_Cb2_X4_0_Xo3(M5_UM5_6_CC8_Cb2_X4_0_NotB, gnd, M5_UM5_6_CC8_Cb2_X4_0_line3);
nand2 M5_UM5_6_CC8_Cb2_X4_0_Xo4(M5_UM5_6_CC8_Cb2_X4_0_line2, M5_UM5_6_CC8_Cb2_X4_0_line3, XCarrybus_0);
inv M5_UM5_6_CC8_Cb2_X4_1_Xo0(M5_UM5_6_CC8_Cy1bus_1, M5_UM5_6_CC8_Cb2_X4_1_NotA);
inv M5_UM5_6_CC8_Cb2_X4_1_Xo1(M5_UM5_6_CC8_Cy2bus_1, M5_UM5_6_CC8_Cb2_X4_1_NotB);
nand2 M5_UM5_6_CC8_Cb2_X4_1_Xo2(M5_UM5_6_CC8_Cb2_X4_1_NotA, M5_UM5_6_CC8_Cy2bus_1, M5_UM5_6_CC8_Cb2_X4_1_line2);
nand2 M5_UM5_6_CC8_Cb2_X4_1_Xo3(M5_UM5_6_CC8_Cb2_X4_1_NotB, M5_UM5_6_CC8_Cy1bus_1, M5_UM5_6_CC8_Cb2_X4_1_line3);
nand2 M5_UM5_6_CC8_Cb2_X4_1_Xo4(M5_UM5_6_CC8_Cb2_X4_1_line2, M5_UM5_6_CC8_Cb2_X4_1_line3, XCarrybus_1);
inv M5_UM5_6_CC8_Cb2_X4_2_Xo0(M5_UM5_6_CC8_Cy1bus_2, M5_UM5_6_CC8_Cb2_X4_2_NotA);
inv M5_UM5_6_CC8_Cb2_X4_2_Xo1(M5_UM5_6_CC8_Cy2bus_2, M5_UM5_6_CC8_Cb2_X4_2_NotB);
nand2 M5_UM5_6_CC8_Cb2_X4_2_Xo2(M5_UM5_6_CC8_Cb2_X4_2_NotA, M5_UM5_6_CC8_Cy2bus_2, M5_UM5_6_CC8_Cb2_X4_2_line2);
nand2 M5_UM5_6_CC8_Cb2_X4_2_Xo3(M5_UM5_6_CC8_Cb2_X4_2_NotB, M5_UM5_6_CC8_Cy1bus_2, M5_UM5_6_CC8_Cb2_X4_2_line3);
nand2 M5_UM5_6_CC8_Cb2_X4_2_Xo4(M5_UM5_6_CC8_Cb2_X4_2_line2, M5_UM5_6_CC8_Cb2_X4_2_line3, XCarrybus_2);
inv M5_UM5_6_CC8_Cb2_X4_3_Xo0(M5_UM5_6_CC8_Cy1bus_3, M5_UM5_6_CC8_Cb2_X4_3_NotA);
inv M5_UM5_6_CC8_Cb2_X4_3_Xo1(M5_UM5_6_CC8_Cy2bus_3, M5_UM5_6_CC8_Cb2_X4_3_NotB);
nand2 M5_UM5_6_CC8_Cb2_X4_3_Xo2(M5_UM5_6_CC8_Cb2_X4_3_NotA, M5_UM5_6_CC8_Cy2bus_3, M5_UM5_6_CC8_Cb2_X4_3_line2);
nand2 M5_UM5_6_CC8_Cb2_X4_3_Xo3(M5_UM5_6_CC8_Cb2_X4_3_NotB, M5_UM5_6_CC8_Cy1bus_3, M5_UM5_6_CC8_Cb2_X4_3_line3);
nand2 M5_UM5_6_CC8_Cb2_X4_3_Xo4(M5_UM5_6_CC8_Cb2_X4_3_line2, M5_UM5_6_CC8_Cb2_X4_3_line3, XCarrybus_3);
and2 M5_UM5_6_CC9_Cb0_Cla4_0_Ao2_0(XPbus_4, M5_UM5_6_LoC0_M, M5_UM5_6_CC9_Cb0_Cla4_0_line0);
or2 M5_UM5_6_CC9_Cb0_Cla4_0_Ao2_1(M5_XGbus_4, M5_UM5_6_CC9_Cb0_Cla4_0_line0, M5_UM5_6_CC9_Cy1bus_1);
and2 M5_UM5_6_CC9_Cb0_Cla4_1_Ao3a_0(XPbus_5, M5_XGbus_4, M5_UM5_6_CC9_Cb0_Cla4_1_line0);
and3 M5_UM5_6_CC9_Cb0_Cla4_1_Ao3a_1(XPbus_5, XPbus_4, M5_UM5_6_LoC0_M, M5_UM5_6_CC9_Cb0_Cla4_1_line1);
or3 M5_UM5_6_CC9_Cb0_Cla4_1_Ao3a_2(M5_XGbus_5, M5_UM5_6_CC9_Cb0_Cla4_1_line0, M5_UM5_6_CC9_Cb0_Cla4_1_line1, M5_UM5_6_CC9_Cy1bus_2);
and2 M5_UM5_6_CC9_Cb0_Cla4_2_Ao4a_0(XPbus_6, M5_XGbus_5, M5_UM5_6_CC9_Cb0_Cla4_2_line0);
and3 M5_UM5_6_CC9_Cb0_Cla4_2_Ao4a_1(XPbus_6, XPbus_5, M5_XGbus_4, M5_UM5_6_CC9_Cb0_Cla4_2_line1);
and4 M5_UM5_6_CC9_Cb0_Cla4_2_Ao4a_2(XPbus_6, XPbus_5, XPbus_4, M5_UM5_6_LoC0_M, M5_UM5_6_CC9_Cb0_Cla4_2_line2);
or4 M5_UM5_6_CC9_Cb0_Cla4_2_Ao4a_3(M5_XGbus_6, M5_UM5_6_CC9_Cb0_Cla4_2_line0, M5_UM5_6_CC9_Cb0_Cla4_2_line1, M5_UM5_6_CC9_Cb0_Cla4_2_line2, M5_UM5_6_CC9_Cy1bus_3);
and2 M5_UM5_6_CC9_Cb1_CP0(XPbus_4, M5_UM5_6_CinPropLo, M5_UM5_6_CC9_Cy2bus_1);
and3 M5_UM5_6_CC9_Cb1_CP1(XPbus_5, XPbus_4, M5_UM5_6_CinPropLo, M5_UM5_6_CC9_Cy2bus_2);
and4 M5_UM5_6_CC9_Cb1_CP2(XPbus_6, XPbus_5, XPbus_4, M5_UM5_6_CinPropLo, M5_UM5_6_CC9_Cy2bus_3);
inv M5_UM5_6_CC9_Cb2_X4_0_Xo0(M5_UM5_6_LoC0_M, M5_UM5_6_CC9_Cb2_X4_0_NotA);
inv M5_UM5_6_CC9_Cb2_X4_0_Xo1(M5_UM5_6_CinPropLo, M5_UM5_6_CC9_Cb2_X4_0_NotB);
nand2 M5_UM5_6_CC9_Cb2_X4_0_Xo2(M5_UM5_6_CC9_Cb2_X4_0_NotA, M5_UM5_6_CinPropLo, M5_UM5_6_CC9_Cb2_X4_0_line2);
nand2 M5_UM5_6_CC9_Cb2_X4_0_Xo3(M5_UM5_6_CC9_Cb2_X4_0_NotB, M5_UM5_6_LoC0_M, M5_UM5_6_CC9_Cb2_X4_0_line3);
nand2 M5_UM5_6_CC9_Cb2_X4_0_Xo4(M5_UM5_6_CC9_Cb2_X4_0_line2, M5_UM5_6_CC9_Cb2_X4_0_line3, XCarrybus_4);
inv M5_UM5_6_CC9_Cb2_X4_1_Xo0(M5_UM5_6_CC9_Cy1bus_1, M5_UM5_6_CC9_Cb2_X4_1_NotA);
inv M5_UM5_6_CC9_Cb2_X4_1_Xo1(M5_UM5_6_CC9_Cy2bus_1, M5_UM5_6_CC9_Cb2_X4_1_NotB);
nand2 M5_UM5_6_CC9_Cb2_X4_1_Xo2(M5_UM5_6_CC9_Cb2_X4_1_NotA, M5_UM5_6_CC9_Cy2bus_1, M5_UM5_6_CC9_Cb2_X4_1_line2);
nand2 M5_UM5_6_CC9_Cb2_X4_1_Xo3(M5_UM5_6_CC9_Cb2_X4_1_NotB, M5_UM5_6_CC9_Cy1bus_1, M5_UM5_6_CC9_Cb2_X4_1_line3);
nand2 M5_UM5_6_CC9_Cb2_X4_1_Xo4(M5_UM5_6_CC9_Cb2_X4_1_line2, M5_UM5_6_CC9_Cb2_X4_1_line3, XCarrybus_5);
inv M5_UM5_6_CC9_Cb2_X4_2_Xo0(M5_UM5_6_CC9_Cy1bus_2, M5_UM5_6_CC9_Cb2_X4_2_NotA);
inv M5_UM5_6_CC9_Cb2_X4_2_Xo1(M5_UM5_6_CC9_Cy2bus_2, M5_UM5_6_CC9_Cb2_X4_2_NotB);
nand2 M5_UM5_6_CC9_Cb2_X4_2_Xo2(M5_UM5_6_CC9_Cb2_X4_2_NotA, M5_UM5_6_CC9_Cy2bus_2, M5_UM5_6_CC9_Cb2_X4_2_line2);
nand2 M5_UM5_6_CC9_Cb2_X4_2_Xo3(M5_UM5_6_CC9_Cb2_X4_2_NotB, M5_UM5_6_CC9_Cy1bus_2, M5_UM5_6_CC9_Cb2_X4_2_line3);
nand2 M5_UM5_6_CC9_Cb2_X4_2_Xo4(M5_UM5_6_CC9_Cb2_X4_2_line2, M5_UM5_6_CC9_Cb2_X4_2_line3, XCarrybus_6);
inv M5_UM5_6_CC9_Cb2_X4_3_Xo0(M5_UM5_6_CC9_Cy1bus_3, M5_UM5_6_CC9_Cb2_X4_3_NotA);
inv M5_UM5_6_CC9_Cb2_X4_3_Xo1(M5_UM5_6_CC9_Cy2bus_3, M5_UM5_6_CC9_Cb2_X4_3_NotB);
nand2 M5_UM5_6_CC9_Cb2_X4_3_Xo2(M5_UM5_6_CC9_Cb2_X4_3_NotA, M5_UM5_6_CC9_Cy2bus_3, M5_UM5_6_CC9_Cb2_X4_3_line2);
nand2 M5_UM5_6_CC9_Cb2_X4_3_Xo3(M5_UM5_6_CC9_Cb2_X4_3_NotB, M5_UM5_6_CC9_Cy1bus_3, M5_UM5_6_CC9_Cb2_X4_3_line3);
nand2 M5_UM5_6_CC9_Cb2_X4_3_Xo4(M5_UM5_6_CC9_Cb2_X4_3_line2, M5_UM5_6_CC9_Cb2_X4_3_line3, XCarrybus_7);
and2 M5_UM5_6_CC10_Ao2_0(M5_UM5_6_LocalC0Lo, M5_UM5_6_PropHi, M5_UM5_6_CC10_line0);
or2 M5_UM5_6_CC10_Ao2_1(M5_UM5_6_LocalC0Hi, M5_UM5_6_CC10_line0, out369);
or2 M5_UM5_6_CC11(M5_UM5_6_CinPropLo, M5_UM5_6_LoC0_M, Carry4);
and2 M5_UM5_6_CC12(M5_UM5_6_CinPropLo, M5_UM5_6_PropHi, M5_UM5_6_line12);
or2 M5_UM5_6_CC13(out369, M5_UM5_6_line12, Cout);
and2 M5_UM5_6_CC14_Ao2_0(M5_UM5_6_LoC0_M, M5_UM5_6_PropHi, M5_UM5_6_CC14_line0);
or2 M5_UM5_6_CC14_Ao2_1(M5_UM5_6_LocalC0Hi, M5_UM5_6_CC14_line0, M5_UM5_6_Cout_M_in0);
inv M5_UM5_6_CC15_Xo0(M5_UM5_6_Cout_M_in0, M5_UM5_6_CC15_NotA);
inv M5_UM5_6_CC15_Xo1(M5_UM5_6_line12, M5_UM5_6_CC15_NotB);
nand2 M5_UM5_6_CC15_Xo2(M5_UM5_6_CC15_NotA, M5_UM5_6_line12, M5_UM5_6_CC15_line2);
nand2 M5_UM5_6_CC15_Xo3(M5_UM5_6_CC15_NotB, M5_UM5_6_Cout_M_in0, M5_UM5_6_CC15_line3);
nand2 M5_UM5_6_CC15_Xo4(M5_UM5_6_CC15_line2, M5_UM5_6_CC15_line3, M5_UM5_6_Ovf_Carry8);
inv M5_UM5_6_CC16_Xo0(M5_UM5_6_Ovf_Carry8, M5_UM5_6_CC16_NotA);
inv M5_UM5_6_CC16_Xo1(XCarrybus_7, M5_UM5_6_CC16_NotB);
nand2 M5_UM5_6_CC16_Xo2(M5_UM5_6_CC16_NotA, XCarrybus_7, M5_UM5_6_CC16_line2);
nand2 M5_UM5_6_CC16_Xo3(M5_UM5_6_CC16_NotB, M5_UM5_6_Ovf_Carry8, M5_UM5_6_CC16_line3);
nand2 M5_UM5_6_CC16_Xo4(M5_UM5_6_CC16_line2, M5_UM5_6_CC16_line3, Overflow);
inv M6_X8_0_X4_0_Xo0(XPbus_0, M6_X8_0_X4_0_NotA);
inv M6_X8_0_X4_0_Xo1(XCarrybus_0, M6_X8_0_X4_0_NotB);
nand2 M6_X8_0_X4_0_Xo2(M6_X8_0_X4_0_NotA, XCarrybus_0, M6_X8_0_X4_0_line2);
nand2 M6_X8_0_X4_0_Xo3(M6_X8_0_X4_0_NotB, XPbus_0, M6_X8_0_X4_0_line3);
nand2 M6_X8_0_X4_0_Xo4(M6_X8_0_X4_0_line2, M6_X8_0_X4_0_line3, Funcbus_0);
inv M6_X8_0_X4_1_Xo0(XPbus_1, M6_X8_0_X4_1_NotA);
inv M6_X8_0_X4_1_Xo1(XCarrybus_1, M6_X8_0_X4_1_NotB);
nand2 M6_X8_0_X4_1_Xo2(M6_X8_0_X4_1_NotA, XCarrybus_1, M6_X8_0_X4_1_line2);
nand2 M6_X8_0_X4_1_Xo3(M6_X8_0_X4_1_NotB, XPbus_1, M6_X8_0_X4_1_line3);
nand2 M6_X8_0_X4_1_Xo4(M6_X8_0_X4_1_line2, M6_X8_0_X4_1_line3, Funcbus_1);
inv M6_X8_0_X4_2_Xo0(XPbus_2, M6_X8_0_X4_2_NotA);
inv M6_X8_0_X4_2_Xo1(XCarrybus_2, M6_X8_0_X4_2_NotB);
nand2 M6_X8_0_X4_2_Xo2(M6_X8_0_X4_2_NotA, XCarrybus_2, M6_X8_0_X4_2_line2);
nand2 M6_X8_0_X4_2_Xo3(M6_X8_0_X4_2_NotB, XPbus_2, M6_X8_0_X4_2_line3);
nand2 M6_X8_0_X4_2_Xo4(M6_X8_0_X4_2_line2, M6_X8_0_X4_2_line3, Funcbus_2);
inv M6_X8_0_X4_3_Xo0(XPbus_3, M6_X8_0_X4_3_NotA);
inv M6_X8_0_X4_3_Xo1(XCarrybus_3, M6_X8_0_X4_3_NotB);
nand2 M6_X8_0_X4_3_Xo2(M6_X8_0_X4_3_NotA, XCarrybus_3, M6_X8_0_X4_3_line2);
nand2 M6_X8_0_X4_3_Xo3(M6_X8_0_X4_3_NotB, XPbus_3, M6_X8_0_X4_3_line3);
nand2 M6_X8_0_X4_3_Xo4(M6_X8_0_X4_3_line2, M6_X8_0_X4_3_line3, Funcbus_3);
inv M6_X8_1_X4_0_Xo0(XPbus_4, M6_X8_1_X4_0_NotA);
inv M6_X8_1_X4_0_Xo1(XCarrybus_4, M6_X8_1_X4_0_NotB);
nand2 M6_X8_1_X4_0_Xo2(M6_X8_1_X4_0_NotA, XCarrybus_4, M6_X8_1_X4_0_line2);
nand2 M6_X8_1_X4_0_Xo3(M6_X8_1_X4_0_NotB, XPbus_4, M6_X8_1_X4_0_line3);
nand2 M6_X8_1_X4_0_Xo4(M6_X8_1_X4_0_line2, M6_X8_1_X4_0_line3, Funcbus_4);
inv M6_X8_1_X4_1_Xo0(XPbus_5, M6_X8_1_X4_1_NotA);
inv M6_X8_1_X4_1_Xo1(XCarrybus_5, M6_X8_1_X4_1_NotB);
nand2 M6_X8_1_X4_1_Xo2(M6_X8_1_X4_1_NotA, XCarrybus_5, M6_X8_1_X4_1_line2);
nand2 M6_X8_1_X4_1_Xo3(M6_X8_1_X4_1_NotB, XPbus_5, M6_X8_1_X4_1_line3);
nand2 M6_X8_1_X4_1_Xo4(M6_X8_1_X4_1_line2, M6_X8_1_X4_1_line3, Funcbus_5);
inv M6_X8_1_X4_2_Xo0(XPbus_6, M6_X8_1_X4_2_NotA);
inv M6_X8_1_X4_2_Xo1(XCarrybus_6, M6_X8_1_X4_2_NotB);
nand2 M6_X8_1_X4_2_Xo2(M6_X8_1_X4_2_NotA, XCarrybus_6, M6_X8_1_X4_2_line2);
nand2 M6_X8_1_X4_2_Xo3(M6_X8_1_X4_2_NotB, XPbus_6, M6_X8_1_X4_2_line3);
nand2 M6_X8_1_X4_2_Xo4(M6_X8_1_X4_2_line2, M6_X8_1_X4_2_line3, Funcbus_6);
inv M6_X8_1_X4_3_Xo0(XPbus_7, M6_X8_1_X4_3_NotA);
inv M6_X8_1_X4_3_Xo1(XCarrybus_7, M6_X8_1_X4_3_NotB);
nand2 M6_X8_1_X4_3_Xo2(M6_X8_1_X4_3_NotA, XCarrybus_7, M6_X8_1_X4_3_line2);
nand2 M6_X8_1_X4_3_Xo3(M6_X8_1_X4_3_NotB, XPbus_7, M6_X8_1_X4_3_line3);
nand2 M6_X8_1_X4_3_Xo4(M6_X8_1_X4_3_line2, M6_X8_1_X4_3_line3, Funcbus_7);
inv M7_UM7_0_Bsd0(Carry4, M7_UM7_0_NotCarry);
inv M7_UM7_0_Bsd1_Xo0(Funcbus_1, M7_UM7_0_Bsd1_NotA);
inv M7_UM7_0_Bsd1_Xo1(M7_UM7_0_NotCarry, M7_UM7_0_Bsd1_NotB);
nand2 M7_UM7_0_Bsd1_Xo2(M7_UM7_0_Bsd1_NotA, M7_UM7_0_NotCarry, M7_UM7_0_Bsd1_line2);
nand2 M7_UM7_0_Bsd1_Xo3(M7_UM7_0_Bsd1_NotB, Funcbus_1, M7_UM7_0_Bsd1_line3);
nand2 M7_UM7_0_Bsd1_Xo4(M7_UM7_0_Bsd1_line2, M7_UM7_0_Bsd1_line3, F_BCDbus_1);
and2 M7_UM7_0_Bsd2(Funcbus_1, M7_UM7_0_NotCarry, M7_UM7_0_line2);
inv M7_UM7_0_Bsd3_Xo0(Funcbus_2, M7_UM7_0_Bsd3_NotA);
inv M7_UM7_0_Bsd3_Xo1(M7_UM7_0_line2, M7_UM7_0_Bsd3_NotB);
nand2 M7_UM7_0_Bsd3_Xo2(M7_UM7_0_Bsd3_NotA, M7_UM7_0_line2, M7_UM7_0_Bsd3_line2);
nand2 M7_UM7_0_Bsd3_Xo3(M7_UM7_0_Bsd3_NotB, Funcbus_2, M7_UM7_0_Bsd3_line3);
nand2 M7_UM7_0_Bsd3_Xo4(M7_UM7_0_Bsd3_line2, M7_UM7_0_Bsd3_line3, F_BCDbus_2);
and4 M7_UM7_0_Bsd4(Funcbus_3, Funcbus_2, Funcbus_1, M7_UM7_0_NotCarry, M7_UM7_0_line4);
and2 M7_UM7_0_Bsd5(Funcbus_3, Carry4, M7_UM7_0_line5);
or2 M7_UM7_0_Bsd6(M7_UM7_0_line4, M7_UM7_0_line5, F_BCDbus_3);
inv M7_UM7_1_Bsd0(Cout, M7_UM7_1_NotCarry);
inv M7_UM7_1_Bsd1_Xo0(Funcbus_5, M7_UM7_1_Bsd1_NotA);
inv M7_UM7_1_Bsd1_Xo1(M7_UM7_1_NotCarry, M7_UM7_1_Bsd1_NotB);
nand2 M7_UM7_1_Bsd1_Xo2(M7_UM7_1_Bsd1_NotA, M7_UM7_1_NotCarry, M7_UM7_1_Bsd1_line2);
nand2 M7_UM7_1_Bsd1_Xo3(M7_UM7_1_Bsd1_NotB, Funcbus_5, M7_UM7_1_Bsd1_line3);
nand2 M7_UM7_1_Bsd1_Xo4(M7_UM7_1_Bsd1_line2, M7_UM7_1_Bsd1_line3, F_BCDbus_5);
and2 M7_UM7_1_Bsd2(Funcbus_5, M7_UM7_1_NotCarry, M7_UM7_1_line2);
inv M7_UM7_1_Bsd3_Xo0(Funcbus_6, M7_UM7_1_Bsd3_NotA);
inv M7_UM7_1_Bsd3_Xo1(M7_UM7_1_line2, M7_UM7_1_Bsd3_NotB);
nand2 M7_UM7_1_Bsd3_Xo2(M7_UM7_1_Bsd3_NotA, M7_UM7_1_line2, M7_UM7_1_Bsd3_line2);
nand2 M7_UM7_1_Bsd3_Xo3(M7_UM7_1_Bsd3_NotB, Funcbus_6, M7_UM7_1_Bsd3_line3);
nand2 M7_UM7_1_Bsd3_Xo4(M7_UM7_1_Bsd3_line2, M7_UM7_1_Bsd3_line3, F_BCDbus_6);
and4 M7_UM7_1_Bsd4(Funcbus_7, Funcbus_6, Funcbus_5, M7_UM7_1_NotCarry, M7_UM7_1_line4);
and2 M7_UM7_1_Bsd5(Funcbus_7, Cout, M7_UM7_1_line5);
or2 M7_UM7_1_Bsd6(M7_UM7_1_line4, M7_UM7_1_line5, F_BCDbus_7);
and2 M8_UM8_0_DCS0(in20, in179, M8_UM8_0_tmp0);
inv M8_UM8_0_DCS1(M8_UM8_0_tmp0, M8_UM8_0_tmp1);
inv M8_UM8_0_DCS2(in20, M8_UM8_0_tmp2);
nand2 M8_UM8_0_DCS3(in20, in200, M8_UM8_0_tmp3);
and2 M8_UM8_0_DCS4(in20, in200, M8_UM8_0_tmp4);
nor2 M8_UM8_0_DCS5(M8_UM8_0_tmp2, in190, M8_UM8_0_tmp5);
and2 M8_UM8_0_DCS6(M8_UM8_0_tmp3, M8_UM8_0_tmp1, M8_UM8_0_tmp6);
and2 M8_UM8_0_DCS7(M8_UM8_0_tmp4, M8_UM8_0_tmp1, M8_UM8_0_tmp7);
or2 M8_UM8_0_DCS8(M8_UM8_0_tmp2, in190, M8_UM8_0_tmp8);
inv M8_UM8_0_DCS9(in200, M8_UM8_0_tmp9);
and2 M8_UM8_0_DCS10(M8_UM8_0_tmp9, M8_UM8_0_tmp0, M8_UM8_0_tmp10);
and2 M8_UM8_0_DCS11(in200, M8_UM8_0_tmp0, M8_UM8_0_tmp11);
and2 M8_UM8_0_DCS13(M8_UM8_0_tmp5, M8_UM8_0_tmp7, M8_ContShift_0);
and2 M8_UM8_0_DCS14(M8_UM8_0_tmp6, M8_UM8_0_tmp8, M8_ContShift_1);
and2 M8_UM8_0_DCS15(M8_UM8_0_tmp8, M8_UM8_0_tmp7, M8_ContShift_2);
and2 M8_UM8_0_DCS16(M8_UM8_0_tmp5, M8_UM8_0_tmp10, M8_ContShift_3);
and2 M8_UM8_0_DCS17(M8_UM8_0_tmp5, M8_UM8_0_tmp11, M8_ContShift_4);
and2 M8_UM8_0_DCS18(M8_UM8_0_tmp8, M8_UM8_0_tmp10, M8_ContShift_5);
and2 M8_UM8_0_DCS19(M8_UM8_0_tmp8, M8_UM8_0_tmp11, M8_ContShift_6);
and2 M8_UM8_0_DCS12(M8_UM8_0_tmp5, M8_UM8_0_tmp6, M8_ContShift_7);
and2 M8_UM8_1_M8_0_M0(in107, M8_ContShift_0, M8_UM8_1_M8_0_t0);
and2 M8_UM8_1_M8_0_M1(in97, M8_ContShift_1, M8_UM8_1_M8_0_t1);
and2 M8_UM8_1_M8_0_M2(in87, M8_ContShift_2, M8_UM8_1_M8_0_t2);
and2 M8_UM8_1_M8_0_M3(in77, M8_ContShift_3, M8_UM8_1_M8_0_t3);
and2 M8_UM8_1_M8_0_M4(in68, M8_ContShift_4, M8_UM8_1_M8_0_t4);
and2 M8_UM8_1_M8_0_M5(in58, M8_ContShift_5, M8_UM8_1_M8_0_t5);
and2 M8_UM8_1_M8_0_M6(in50, M8_ContShift_6, M8_UM8_1_M8_0_t6);
and2 M8_UM8_1_M8_0_M7(in159, M8_ContShift_7, M8_UM8_1_M8_0_t7);
or8 M8_UM8_1_M8_0_M8(M8_UM8_1_M8_0_t0, M8_UM8_1_M8_0_t1, M8_UM8_1_M8_0_t2, M8_UM8_1_M8_0_t3, M8_UM8_1_M8_0_t4, M8_UM8_1_M8_0_t5, M8_UM8_1_M8_0_t6, M8_UM8_1_M8_0_t7, M8_ShiftQout_0);
and2 M8_UM8_1_M8_1_M0(in97, M8_ContShift_0, M8_UM8_1_M8_1_t0);
and2 M8_UM8_1_M8_1_M1(in87, M8_ContShift_1, M8_UM8_1_M8_1_t1);
and2 M8_UM8_1_M8_1_M2(in77, M8_ContShift_2, M8_UM8_1_M8_1_t2);
and2 M8_UM8_1_M8_1_M3(in68, M8_ContShift_3, M8_UM8_1_M8_1_t3);
and2 M8_UM8_1_M8_1_M4(in58, M8_ContShift_4, M8_UM8_1_M8_1_t4);
and2 M8_UM8_1_M8_1_M5(in50, M8_ContShift_5, M8_UM8_1_M8_1_t5);
and2 M8_UM8_1_M8_1_M6(in159, M8_ContShift_6, M8_UM8_1_M8_1_t6);
and2 M8_UM8_1_M8_1_M7(in150, M8_ContShift_7, M8_UM8_1_M8_1_t7);
or8 M8_UM8_1_M8_1_M8(M8_UM8_1_M8_1_t0, M8_UM8_1_M8_1_t1, M8_UM8_1_M8_1_t2, M8_UM8_1_M8_1_t3, M8_UM8_1_M8_1_t4, M8_UM8_1_M8_1_t5, M8_UM8_1_M8_1_t6, M8_UM8_1_M8_1_t7, M8_ShiftQout_1);
and2 M8_UM8_1_M8_2_M0(in87, M8_ContShift_0, M8_UM8_1_M8_2_t0);
and2 M8_UM8_1_M8_2_M1(in77, M8_ContShift_1, M8_UM8_1_M8_2_t1);
and2 M8_UM8_1_M8_2_M2(in68, M8_ContShift_2, M8_UM8_1_M8_2_t2);
and2 M8_UM8_1_M8_2_M3(in58, M8_ContShift_3, M8_UM8_1_M8_2_t3);
and2 M8_UM8_1_M8_2_M4(in50, M8_ContShift_4, M8_UM8_1_M8_2_t4);
and2 M8_UM8_1_M8_2_M5(in159, M8_ContShift_5, M8_UM8_1_M8_2_t5);
and2 M8_UM8_1_M8_2_M6(in150, M8_ContShift_6, M8_UM8_1_M8_2_t6);
and2 M8_UM8_1_M8_2_M7(in143, M8_ContShift_7, M8_UM8_1_M8_2_t7);
or8 M8_UM8_1_M8_2_M8(M8_UM8_1_M8_2_t0, M8_UM8_1_M8_2_t1, M8_UM8_1_M8_2_t2, M8_UM8_1_M8_2_t3, M8_UM8_1_M8_2_t4, M8_UM8_1_M8_2_t5, M8_UM8_1_M8_2_t6, M8_UM8_1_M8_2_t7, M8_ShiftQout_2);
and2 M8_UM8_1_M8_3_M0(in77, M8_ContShift_0, M8_UM8_1_M8_3_t0);
and2 M8_UM8_1_M8_3_M1(in68, M8_ContShift_1, M8_UM8_1_M8_3_t1);
and2 M8_UM8_1_M8_3_M2(in58, M8_ContShift_2, M8_UM8_1_M8_3_t2);
and2 M8_UM8_1_M8_3_M3(in50, M8_ContShift_3, M8_UM8_1_M8_3_t3);
and2 M8_UM8_1_M8_3_M4(in159, M8_ContShift_4, M8_UM8_1_M8_3_t4);
and2 M8_UM8_1_M8_3_M5(in150, M8_ContShift_5, M8_UM8_1_M8_3_t5);
and2 M8_UM8_1_M8_3_M6(in143, M8_ContShift_6, M8_UM8_1_M8_3_t6);
and2 M8_UM8_1_M8_3_M7(in137, M8_ContShift_7, M8_UM8_1_M8_3_t7);
or8 M8_UM8_1_M8_3_M8(M8_UM8_1_M8_3_t0, M8_UM8_1_M8_3_t1, M8_UM8_1_M8_3_t2, M8_UM8_1_M8_3_t3, M8_UM8_1_M8_3_t4, M8_UM8_1_M8_3_t5, M8_UM8_1_M8_3_t6, M8_UM8_1_M8_3_t7, M8_ShiftQout_3);
and2 M8_UM8_1_M8_4_M0(in68, M8_ContShift_0, M8_UM8_1_M8_4_t0);
and2 M8_UM8_1_M8_4_M1(in58, M8_ContShift_1, M8_UM8_1_M8_4_t1);
and2 M8_UM8_1_M8_4_M2(in50, M8_ContShift_2, M8_UM8_1_M8_4_t2);
and2 M8_UM8_1_M8_4_M3(in159, M8_ContShift_3, M8_UM8_1_M8_4_t3);
and2 M8_UM8_1_M8_4_M4(in150, M8_ContShift_4, M8_UM8_1_M8_4_t4);
and2 M8_UM8_1_M8_4_M5(in143, M8_ContShift_5, M8_UM8_1_M8_4_t5);
and2 M8_UM8_1_M8_4_M6(in137, M8_ContShift_6, M8_UM8_1_M8_4_t6);
and2 M8_UM8_1_M8_4_M7(in132, M8_ContShift_7, M8_UM8_1_M8_4_t7);
or8 M8_UM8_1_M8_4_M8(M8_UM8_1_M8_4_t0, M8_UM8_1_M8_4_t1, M8_UM8_1_M8_4_t2, M8_UM8_1_M8_4_t3, M8_UM8_1_M8_4_t4, M8_UM8_1_M8_4_t5, M8_UM8_1_M8_4_t6, M8_UM8_1_M8_4_t7, M8_ShiftQout_4);
and2 M8_UM8_1_M8_5_M0(in58, M8_ContShift_0, M8_UM8_1_M8_5_t0);
and2 M8_UM8_1_M8_5_M1(in50, M8_ContShift_1, M8_UM8_1_M8_5_t1);
and2 M8_UM8_1_M8_5_M2(in159, M8_ContShift_2, M8_UM8_1_M8_5_t2);
and2 M8_UM8_1_M8_5_M3(in150, M8_ContShift_3, M8_UM8_1_M8_5_t3);
and2 M8_UM8_1_M8_5_M4(in143, M8_ContShift_4, M8_UM8_1_M8_5_t4);
and2 M8_UM8_1_M8_5_M5(in137, M8_ContShift_5, M8_UM8_1_M8_5_t5);
and2 M8_UM8_1_M8_5_M6(in132, M8_ContShift_6, M8_UM8_1_M8_5_t6);
and2 M8_UM8_1_M8_5_M7(in128, M8_ContShift_7, M8_UM8_1_M8_5_t7);
or8 M8_UM8_1_M8_5_M8(M8_UM8_1_M8_5_t0, M8_UM8_1_M8_5_t1, M8_UM8_1_M8_5_t2, M8_UM8_1_M8_5_t3, M8_UM8_1_M8_5_t4, M8_UM8_1_M8_5_t5, M8_UM8_1_M8_5_t6, M8_UM8_1_M8_5_t7, M8_ShiftQout_5);
and2 M8_UM8_1_M8_6_M0(in50, M8_ContShift_0, M8_UM8_1_M8_6_t0);
and2 M8_UM8_1_M8_6_M1(in159, M8_ContShift_1, M8_UM8_1_M8_6_t1);
and2 M8_UM8_1_M8_6_M2(in150, M8_ContShift_2, M8_UM8_1_M8_6_t2);
and2 M8_UM8_1_M8_6_M3(in143, M8_ContShift_3, M8_UM8_1_M8_6_t3);
and2 M8_UM8_1_M8_6_M4(in137, M8_ContShift_4, M8_UM8_1_M8_6_t4);
and2 M8_UM8_1_M8_6_M5(in132, M8_ContShift_5, M8_UM8_1_M8_6_t5);
and2 M8_UM8_1_M8_6_M6(in128, M8_ContShift_6, M8_UM8_1_M8_6_t6);
and2 M8_UM8_1_M8_6_M7(in125, M8_ContShift_7, M8_UM8_1_M8_6_t7);
or8 M8_UM8_1_M8_6_M8(M8_UM8_1_M8_6_t0, M8_UM8_1_M8_6_t1, M8_UM8_1_M8_6_t2, M8_UM8_1_M8_6_t3, M8_UM8_1_M8_6_t4, M8_UM8_1_M8_6_t5, M8_UM8_1_M8_6_t6, M8_UM8_1_M8_6_t7, M8_ShiftQout_6);
and2 M8_UM8_1_M8_7_M0(in159, M8_ContShift_0, M8_UM8_1_M8_7_t0);
and2 M8_UM8_1_M8_7_M1(in150, M8_ContShift_1, M8_UM8_1_M8_7_t1);
and2 M8_UM8_1_M8_7_M2(in143, M8_ContShift_2, M8_UM8_1_M8_7_t2);
and2 M8_UM8_1_M8_7_M3(in137, M8_ContShift_3, M8_UM8_1_M8_7_t3);
and2 M8_UM8_1_M8_7_M4(in132, M8_ContShift_4, M8_UM8_1_M8_7_t4);
and2 M8_UM8_1_M8_7_M5(in128, M8_ContShift_5, M8_UM8_1_M8_7_t5);
and2 M8_UM8_1_M8_7_M6(in125, M8_ContShift_6, M8_UM8_1_M8_7_t6);
and2 M8_UM8_1_M8_7_M7(in124, M8_ContShift_7, M8_UM8_1_M8_7_t7);
or8 M8_UM8_1_M8_7_M8(M8_UM8_1_M8_7_t0, M8_UM8_1_M8_7_t1, M8_UM8_1_M8_7_t2, M8_UM8_1_M8_7_t3, M8_UM8_1_M8_7_t4, M8_UM8_1_M8_7_t5, M8_UM8_1_M8_7_t6, M8_UM8_1_M8_7_t7, M8_ShiftQout_7);
and2 M8_UM8_2_M8_0_M0(in283, M8_ContShift_0, M8_UM8_2_M8_0_t0);
and2 M8_UM8_2_M8_0_M1(in294, M8_ContShift_1, M8_UM8_2_M8_0_t1);
and2 M8_UM8_2_M8_0_M2(in303, M8_ContShift_2, M8_UM8_2_M8_0_t2);
and2 M8_UM8_2_M8_0_M3(in311, M8_ContShift_3, M8_UM8_2_M8_0_t3);
and2 M8_UM8_2_M8_0_M4(in317, M8_ContShift_4, M8_UM8_2_M8_0_t4);
and2 M8_UM8_2_M8_0_M5(in322, M8_ContShift_5, M8_UM8_2_M8_0_t5);
and2 M8_UM8_2_M8_0_M6(in326, M8_ContShift_6, M8_UM8_2_M8_0_t6);
and2 M8_UM8_2_M8_0_M7(in329, M8_ContShift_7, M8_UM8_2_M8_0_t7);
or8 M8_UM8_2_M8_0_M8(M8_UM8_2_M8_0_t0, M8_UM8_2_M8_0_t1, M8_UM8_2_M8_0_t2, M8_UM8_2_M8_0_t3, M8_UM8_2_M8_0_t4, M8_UM8_2_M8_0_t5, M8_UM8_2_M8_0_t6, M8_UM8_2_M8_0_t7, M8_ShiftRout_0);
and2 M8_UM8_2_M8_1_M0(in116, M8_ContShift_0, M8_UM8_2_M8_1_t0);
and2 M8_UM8_2_M8_1_M1(in283, M8_ContShift_1, M8_UM8_2_M8_1_t1);
and2 M8_UM8_2_M8_1_M2(in294, M8_ContShift_2, M8_UM8_2_M8_1_t2);
and2 M8_UM8_2_M8_1_M3(in303, M8_ContShift_3, M8_UM8_2_M8_1_t3);
and2 M8_UM8_2_M8_1_M4(in311, M8_ContShift_4, M8_UM8_2_M8_1_t4);
and2 M8_UM8_2_M8_1_M5(in317, M8_ContShift_5, M8_UM8_2_M8_1_t5);
and2 M8_UM8_2_M8_1_M6(in322, M8_ContShift_6, M8_UM8_2_M8_1_t6);
and2 M8_UM8_2_M8_1_M7(in326, M8_ContShift_7, M8_UM8_2_M8_1_t7);
or8 M8_UM8_2_M8_1_M8(M8_UM8_2_M8_1_t0, M8_UM8_2_M8_1_t1, M8_UM8_2_M8_1_t2, M8_UM8_2_M8_1_t3, M8_UM8_2_M8_1_t4, M8_UM8_2_M8_1_t5, M8_UM8_2_M8_1_t6, M8_UM8_2_M8_1_t7, M8_ShiftRout_1);
and2 M8_UM8_2_M8_2_M0(in107, M8_ContShift_0, M8_UM8_2_M8_2_t0);
and2 M8_UM8_2_M8_2_M1(in116, M8_ContShift_1, M8_UM8_2_M8_2_t1);
and2 M8_UM8_2_M8_2_M2(in283, M8_ContShift_2, M8_UM8_2_M8_2_t2);
and2 M8_UM8_2_M8_2_M3(in294, M8_ContShift_3, M8_UM8_2_M8_2_t3);
and2 M8_UM8_2_M8_2_M4(in303, M8_ContShift_4, M8_UM8_2_M8_2_t4);
and2 M8_UM8_2_M8_2_M5(in311, M8_ContShift_5, M8_UM8_2_M8_2_t5);
and2 M8_UM8_2_M8_2_M6(in317, M8_ContShift_6, M8_UM8_2_M8_2_t6);
and2 M8_UM8_2_M8_2_M7(in322, M8_ContShift_7, M8_UM8_2_M8_2_t7);
or8 M8_UM8_2_M8_2_M8(M8_UM8_2_M8_2_t0, M8_UM8_2_M8_2_t1, M8_UM8_2_M8_2_t2, M8_UM8_2_M8_2_t3, M8_UM8_2_M8_2_t4, M8_UM8_2_M8_2_t5, M8_UM8_2_M8_2_t6, M8_UM8_2_M8_2_t7, M8_ShiftRout_2);
and2 M8_UM8_2_M8_3_M0(in97, M8_ContShift_0, M8_UM8_2_M8_3_t0);
and2 M8_UM8_2_M8_3_M1(in107, M8_ContShift_1, M8_UM8_2_M8_3_t1);
and2 M8_UM8_2_M8_3_M2(in116, M8_ContShift_2, M8_UM8_2_M8_3_t2);
and2 M8_UM8_2_M8_3_M3(in283, M8_ContShift_3, M8_UM8_2_M8_3_t3);
and2 M8_UM8_2_M8_3_M4(in294, M8_ContShift_4, M8_UM8_2_M8_3_t4);
and2 M8_UM8_2_M8_3_M5(in303, M8_ContShift_5, M8_UM8_2_M8_3_t5);
and2 M8_UM8_2_M8_3_M6(in311, M8_ContShift_6, M8_UM8_2_M8_3_t6);
and2 M8_UM8_2_M8_3_M7(in317, M8_ContShift_7, M8_UM8_2_M8_3_t7);
or8 M8_UM8_2_M8_3_M8(M8_UM8_2_M8_3_t0, M8_UM8_2_M8_3_t1, M8_UM8_2_M8_3_t2, M8_UM8_2_M8_3_t3, M8_UM8_2_M8_3_t4, M8_UM8_2_M8_3_t5, M8_UM8_2_M8_3_t6, M8_UM8_2_M8_3_t7, M8_ShiftRout_3);
and2 M8_UM8_2_M8_4_M0(in87, M8_ContShift_0, M8_UM8_2_M8_4_t0);
and2 M8_UM8_2_M8_4_M1(in97, M8_ContShift_1, M8_UM8_2_M8_4_t1);
and2 M8_UM8_2_M8_4_M2(in107, M8_ContShift_2, M8_UM8_2_M8_4_t2);
and2 M8_UM8_2_M8_4_M3(in116, M8_ContShift_3, M8_UM8_2_M8_4_t3);
and2 M8_UM8_2_M8_4_M4(in283, M8_ContShift_4, M8_UM8_2_M8_4_t4);
and2 M8_UM8_2_M8_4_M5(in294, M8_ContShift_5, M8_UM8_2_M8_4_t5);
and2 M8_UM8_2_M8_4_M6(in303, M8_ContShift_6, M8_UM8_2_M8_4_t6);
and2 M8_UM8_2_M8_4_M7(in311, M8_ContShift_7, M8_UM8_2_M8_4_t7);
or8 M8_UM8_2_M8_4_M8(M8_UM8_2_M8_4_t0, M8_UM8_2_M8_4_t1, M8_UM8_2_M8_4_t2, M8_UM8_2_M8_4_t3, M8_UM8_2_M8_4_t4, M8_UM8_2_M8_4_t5, M8_UM8_2_M8_4_t6, M8_UM8_2_M8_4_t7, M8_ShiftRout_4);
and2 M8_UM8_2_M8_5_M0(in77, M8_ContShift_0, M8_UM8_2_M8_5_t0);
and2 M8_UM8_2_M8_5_M1(in87, M8_ContShift_1, M8_UM8_2_M8_5_t1);
and2 M8_UM8_2_M8_5_M2(in97, M8_ContShift_2, M8_UM8_2_M8_5_t2);
and2 M8_UM8_2_M8_5_M3(in107, M8_ContShift_3, M8_UM8_2_M8_5_t3);
and2 M8_UM8_2_M8_5_M4(in116, M8_ContShift_4, M8_UM8_2_M8_5_t4);
and2 M8_UM8_2_M8_5_M5(in283, M8_ContShift_5, M8_UM8_2_M8_5_t5);
and2 M8_UM8_2_M8_5_M6(in294, M8_ContShift_6, M8_UM8_2_M8_5_t6);
and2 M8_UM8_2_M8_5_M7(in303, M8_ContShift_7, M8_UM8_2_M8_5_t7);
or8 M8_UM8_2_M8_5_M8(M8_UM8_2_M8_5_t0, M8_UM8_2_M8_5_t1, M8_UM8_2_M8_5_t2, M8_UM8_2_M8_5_t3, M8_UM8_2_M8_5_t4, M8_UM8_2_M8_5_t5, M8_UM8_2_M8_5_t6, M8_UM8_2_M8_5_t7, M8_ShiftRout_5);
and2 M8_UM8_2_M8_6_M0(in68, M8_ContShift_0, M8_UM8_2_M8_6_t0);
and2 M8_UM8_2_M8_6_M1(in77, M8_ContShift_1, M8_UM8_2_M8_6_t1);
and2 M8_UM8_2_M8_6_M2(in87, M8_ContShift_2, M8_UM8_2_M8_6_t2);
and2 M8_UM8_2_M8_6_M3(in97, M8_ContShift_3, M8_UM8_2_M8_6_t3);
and2 M8_UM8_2_M8_6_M4(in107, M8_ContShift_4, M8_UM8_2_M8_6_t4);
and2 M8_UM8_2_M8_6_M5(in116, M8_ContShift_5, M8_UM8_2_M8_6_t5);
and2 M8_UM8_2_M8_6_M6(in283, M8_ContShift_6, M8_UM8_2_M8_6_t6);
and2 M8_UM8_2_M8_6_M7(in294, M8_ContShift_7, M8_UM8_2_M8_6_t7);
or8 M8_UM8_2_M8_6_M8(M8_UM8_2_M8_6_t0, M8_UM8_2_M8_6_t1, M8_UM8_2_M8_6_t2, M8_UM8_2_M8_6_t3, M8_UM8_2_M8_6_t4, M8_UM8_2_M8_6_t5, M8_UM8_2_M8_6_t6, M8_UM8_2_M8_6_t7, M8_ShiftRout_6);
and2 M8_UM8_2_M8_7_M0(in58, M8_ContShift_0, M8_UM8_2_M8_7_t0);
and2 M8_UM8_2_M8_7_M1(in68, M8_ContShift_1, M8_UM8_2_M8_7_t1);
and2 M8_UM8_2_M8_7_M2(in77, M8_ContShift_2, M8_UM8_2_M8_7_t2);
and2 M8_UM8_2_M8_7_M3(in87, M8_ContShift_3, M8_UM8_2_M8_7_t3);
and2 M8_UM8_2_M8_7_M4(in97, M8_ContShift_4, M8_UM8_2_M8_7_t4);
and2 M8_UM8_2_M8_7_M5(in107, M8_ContShift_5, M8_UM8_2_M8_7_t5);
and2 M8_UM8_2_M8_7_M6(in116, M8_ContShift_6, M8_UM8_2_M8_7_t6);
and2 M8_UM8_2_M8_7_M7(in283, M8_ContShift_7, M8_UM8_2_M8_7_t7);
or8 M8_UM8_2_M8_7_M8(M8_UM8_2_M8_7_t0, M8_UM8_2_M8_7_t1, M8_UM8_2_M8_7_t2, M8_UM8_2_M8_7_t3, M8_UM8_2_M8_7_t4, M8_UM8_2_M8_7_t5, M8_UM8_2_M8_7_t6, M8_UM8_2_M8_7_t7, M8_ShiftRout_7);
inv M8_UM8_3_Mux2_0(in33, M8_UM8_3_Not_ContIn);
and2 M8_UM8_3_Mux2_1(M8_ShiftQout_0, M8_UM8_3_Not_ContIn, M8_UM8_3_line1);
and2 M8_UM8_3_Mux2_2(M8_ShiftRout_0, in33, M8_UM8_3_line2);
or2 M8_UM8_3_Mux2_3(M8_UM8_3_line1, M8_UM8_3_line2, Shiftbus_0);
inv M8_UM8_4_Mux2_0(in33, M8_UM8_4_Not_ContIn);
and2 M8_UM8_4_Mux2_1(M8_ShiftQout_1, M8_UM8_4_Not_ContIn, M8_UM8_4_line1);
and2 M8_UM8_4_Mux2_2(M8_ShiftRout_1, in33, M8_UM8_4_line2);
or2 M8_UM8_4_Mux2_3(M8_UM8_4_line1, M8_UM8_4_line2, Shiftbus_1);
inv M8_UM8_5_Mux2_0(in33, M8_UM8_5_Not_ContIn);
and2 M8_UM8_5_Mux2_1(M8_ShiftQout_2, M8_UM8_5_Not_ContIn, M8_UM8_5_line1);
and2 M8_UM8_5_Mux2_2(M8_ShiftRout_2, in33, M8_UM8_5_line2);
or2 M8_UM8_5_Mux2_3(M8_UM8_5_line1, M8_UM8_5_line2, Shiftbus_2);
inv M8_UM8_6_Mux2_0(in33, M8_UM8_6_Not_ContIn);
and2 M8_UM8_6_Mux2_1(M8_ShiftQout_3, M8_UM8_6_Not_ContIn, M8_UM8_6_line1);
and2 M8_UM8_6_Mux2_2(M8_ShiftRout_3, in33, M8_UM8_6_line2);
or2 M8_UM8_6_Mux2_3(M8_UM8_6_line1, M8_UM8_6_line2, Shiftbus_3);
inv M8_UM8_7_Mux2_0(in33, M8_UM8_7_Not_ContIn);
and2 M8_UM8_7_Mux2_1(M8_ShiftQout_4, M8_UM8_7_Not_ContIn, M8_UM8_7_line1);
and2 M8_UM8_7_Mux2_2(M8_ShiftRout_4, in33, M8_UM8_7_line2);
or2 M8_UM8_7_Mux2_3(M8_UM8_7_line1, M8_UM8_7_line2, Shiftbus_4);
inv M8_UM8_8_Mux2_0(in33, M8_UM8_8_Not_ContIn);
and2 M8_UM8_8_Mux2_1(M8_ShiftQout_5, M8_UM8_8_Not_ContIn, M8_UM8_8_line1);
and2 M8_UM8_8_Mux2_2(M8_ShiftRout_5, in33, M8_UM8_8_line2);
or2 M8_UM8_8_Mux2_3(M8_UM8_8_line1, M8_UM8_8_line2, Shiftbus_5);
inv M8_UM8_9_Mux2_0(in33, M8_UM8_9_Not_ContIn);
and2 M8_UM8_9_Mux2_1(M8_ShiftQout_6, M8_UM8_9_Not_ContIn, M8_UM8_9_line1);
and2 M8_UM8_9_Mux2_2(M8_ShiftRout_6, in33, M8_UM8_9_line2);
or2 M8_UM8_9_Mux2_3(M8_UM8_9_line1, M8_UM8_9_line2, Shiftbus_6);
inv M8_UM8_10_Mux2_0(in33, M8_UM8_10_Not_ContIn);
and2 M8_UM8_10_Mux2_1(M8_ShiftQout_7, M8_UM8_10_Not_ContIn, M8_UM8_10_line1);
and2 M8_UM8_10_Mux2_2(M8_ShiftRout_7, in33, M8_UM8_10_line2);
or2 M8_UM8_10_Mux2_3(M8_UM8_10_line1, M8_UM8_10_line2, M8_Sbus7_0);
inv M8_UM8_11_Mux2_0(in41, M8_UM8_11_Not_ContIn);
and2 M8_UM8_11_Mux2_1(M8_Sbus7_0, M8_UM8_11_Not_ContIn, M8_UM8_11_line1);
and2 M8_UM8_11_Mux2_2(in50, in41, M8_UM8_11_line2);
or2 M8_UM8_11_Mux2_3(M8_UM8_11_line1, M8_UM8_11_line2, Shiftbus_7);
inv M9_UM9_0_BM0_Inv8_0_Inv4_0(in116, M9_UM9_0_NotAbus_0);
inv M9_UM9_0_BM0_Inv8_0_Inv4_1(in107, M9_UM9_0_NotAbus_1);
inv M9_UM9_0_BM0_Inv8_0_Inv4_2(in97, M9_UM9_0_NotAbus_2);
inv M9_UM9_0_BM0_Inv8_0_Inv4_3(in87, M9_UM9_0_NotAbus_3);
inv M9_UM9_0_BM0_Inv8_1_Inv4_0(in77, M9_UM9_0_NotAbus_4);
inv M9_UM9_0_BM0_Inv8_1_Inv4_1(in68, M9_UM9_0_NotAbus_5);
inv M9_UM9_0_BM0_Inv8_1_Inv4_2(in58, M9_UM9_0_NotAbus_6);
inv M9_UM9_0_BM0_Inv8_1_Inv4_3(in50, M9_UM9_0_NotAbus_7);
nand2 M9_UM9_0_BM1(M9_UM9_0_NotAbus_6, M9_UM9_0_NotAbus_5, M9_UM9_0_NotA6_5);
and2 M9_UM9_0_BM2(in50, M9_UM9_0_NotA6_5, M9_UM9_0_T1_0_0);
inv M9_UM9_0_BM3_Xo0(M9_UM9_0_NotAbus_4, M9_UM9_0_BM3_NotA);
inv M9_UM9_0_BM3_Xo1(M9_UM9_0_NotAbus_5, M9_UM9_0_BM3_NotB);
nand2 M9_UM9_0_BM3_Xo2(M9_UM9_0_BM3_NotA, M9_UM9_0_NotAbus_5, M9_UM9_0_BM3_line2);
nand2 M9_UM9_0_BM3_Xo3(M9_UM9_0_BM3_NotB, M9_UM9_0_NotAbus_4, M9_UM9_0_BM3_line3);
nand2 M9_UM9_0_BM3_Xo4(M9_UM9_0_BM3_line2, M9_UM9_0_BM3_line3, M9_UM9_0_XA5_4);
inv M9_UM9_0_BM4_Xo0(M9_UM9_0_NotAbus_6, M9_UM9_0_BM4_NotA);
inv M9_UM9_0_BM4_Xo1(in50, M9_UM9_0_BM4_NotB);
nand2 M9_UM9_0_BM4_Xo2(M9_UM9_0_BM4_NotA, in50, M9_UM9_0_BM4_line2);
nand2 M9_UM9_0_BM4_Xo3(M9_UM9_0_BM4_NotB, M9_UM9_0_NotAbus_6, M9_UM9_0_BM4_line3);
nand2 M9_UM9_0_BM4_Xo4(M9_UM9_0_BM4_line2, M9_UM9_0_BM4_line3, M9_UM9_0_NotXA7_6);
inv M9_UM9_0_BM5_Xo0(M9_UM9_0_XA5_4, M9_UM9_0_BM5_NotA);
inv M9_UM9_0_BM5_Xo1(M9_UM9_0_NotXA7_6, M9_UM9_0_BM5_NotB);
nand2 M9_UM9_0_BM5_Xo2(M9_UM9_0_BM5_NotA, M9_UM9_0_NotXA7_6, M9_UM9_0_BM5_line2);
nand2 M9_UM9_0_BM5_Xo3(M9_UM9_0_BM5_NotB, M9_UM9_0_XA5_4, M9_UM9_0_BM5_line3);
nand2 M9_UM9_0_BM5_Xo4(M9_UM9_0_BM5_line2, M9_UM9_0_BM5_line3, M9_UM9_0_T1_0_1);
inv M9_UM9_0_BM6_Mux2_0(in45, M9_UM9_0_BM6_Not_ContIn);
and2 M9_UM9_0_BM6_Mux2_1(M9_UM9_0_T1_0_0, M9_UM9_0_BM6_Not_ContIn, M9_UM9_0_BM6_line1);
and2 M9_UM9_0_BM6_Mux2_2(M9_UM9_0_T1_0_1, in45, M9_UM9_0_BM6_line2);
or2 M9_UM9_0_BM6_Mux2_3(M9_UM9_0_BM6_line1, M9_UM9_0_BM6_line2, M9_temp1bus_0);
and3 M9_UM9_0_BM7(M9_UM9_0_NotAbus_3, M9_UM9_0_NotAbus_2, M9_UM9_0_NotAbus_1, M9_UM9_0_NotA3_1);
and2 M9_UM9_0_BM8(M9_UM9_0_NotAbus_0, M9_UM9_0_NotA3_1, M9_UM9_0_NotA3_0);
nand2 M9_UM9_0_BM9(in77, in68, M9_UM9_0_NdA5_4);
and4 M9_UM9_0_BM10(M9_UM9_0_NotA3_0, M9_UM9_0_NdA5_4, M9_UM9_0_NotAbus_7, in58, M9_UM9_0_T1_1_0);
inv M9_UM9_0_BM11_Xo0(in244, M9_UM9_0_BM11_NotA);
inv M9_UM9_0_BM11_Xo1(in238, M9_UM9_0_BM11_NotB);
nand2 M9_UM9_0_BM11_Xo2(M9_UM9_0_BM11_NotA, in238, M9_UM9_0_BM11_line2);
nand2 M9_UM9_0_BM11_Xo3(M9_UM9_0_BM11_NotB, in244, M9_UM9_0_BM11_line3);
nand2 M9_UM9_0_BM11_Xo4(M9_UM9_0_BM11_line2, M9_UM9_0_BM11_line3, M9_UM9_0_XB5_4);
inv M9_UM9_0_BM12_Xo0(in226, M9_UM9_0_BM12_NotA);
inv M9_UM9_0_BM12_Xo1(in232, M9_UM9_0_BM12_NotB);
nand2 M9_UM9_0_BM12_Xo2(M9_UM9_0_BM12_NotA, in232, M9_UM9_0_BM12_line2);
nand2 M9_UM9_0_BM12_Xo3(M9_UM9_0_BM12_NotB, in226, M9_UM9_0_BM12_line3);
nand2 M9_UM9_0_BM12_Xo4(M9_UM9_0_BM12_line2, M9_UM9_0_BM12_line3, M9_UM9_0_XB7_6);
inv M9_UM9_0_BM13_Xo0(M9_UM9_0_XB5_4, M9_UM9_0_BM13_NotA);
inv M9_UM9_0_BM13_Xo1(M9_UM9_0_XB7_6, M9_UM9_0_BM13_NotB);
nand2 M9_UM9_0_BM13_Xo2(M9_UM9_0_BM13_NotA, M9_UM9_0_XB7_6, M9_UM9_0_BM13_line2);
nand2 M9_UM9_0_BM13_Xo3(M9_UM9_0_BM13_NotB, M9_UM9_0_XB5_4, M9_UM9_0_BM13_line3);
nand2 M9_UM9_0_BM13_Xo4(M9_UM9_0_BM13_line2, M9_UM9_0_BM13_line3, M9_UM9_0_XB7_4);
inv M9_UM9_0_BM14(M9_UM9_0_XB7_4, M9_UM9_0_T1_1_1);
inv M9_UM9_0_BM15_Mux2_0(in45, M9_UM9_0_BM15_Not_ContIn);
and2 M9_UM9_0_BM15_Mux2_1(M9_UM9_0_T1_1_0, M9_UM9_0_BM15_Not_ContIn, M9_UM9_0_BM15_line1);
and2 M9_UM9_0_BM15_Mux2_2(M9_UM9_0_T1_1_1, in45, M9_UM9_0_BM15_line2);
or2 M9_UM9_0_BM15_Mux2_3(M9_UM9_0_BM15_line1, M9_UM9_0_BM15_line2, M9_temp1bus_1);
inv M9_UM9_0_BM16_Xo0(M9_UM9_0_NotAbus_0, M9_UM9_0_BM16_NotA);
inv M9_UM9_0_BM16_Xo1(M9_UM9_0_NotAbus_1, M9_UM9_0_BM16_NotB);
nand2 M9_UM9_0_BM16_Xo2(M9_UM9_0_BM16_NotA, M9_UM9_0_NotAbus_1, M9_UM9_0_BM16_line2);
nand2 M9_UM9_0_BM16_Xo3(M9_UM9_0_BM16_NotB, M9_UM9_0_NotAbus_0, M9_UM9_0_BM16_line3);
nand2 M9_UM9_0_BM16_Xo4(M9_UM9_0_BM16_line2, M9_UM9_0_BM16_line3, M9_UM9_0_XA1_0);
inv M9_UM9_0_BM17_Xo0(M9_UM9_0_NotAbus_2, M9_UM9_0_BM17_NotA);
inv M9_UM9_0_BM17_Xo1(M9_UM9_0_NotAbus_3, M9_UM9_0_BM17_NotB);
nand2 M9_UM9_0_BM17_Xo2(M9_UM9_0_BM17_NotA, M9_UM9_0_NotAbus_3, M9_UM9_0_BM17_line2);
nand2 M9_UM9_0_BM17_Xo3(M9_UM9_0_BM17_NotB, M9_UM9_0_NotAbus_2, M9_UM9_0_BM17_line3);
nand2 M9_UM9_0_BM17_Xo4(M9_UM9_0_BM17_line2, M9_UM9_0_BM17_line3, M9_UM9_0_XA3_2);
inv M9_UM9_0_BM18_Xo0(M9_UM9_0_XA1_0, M9_UM9_0_BM18_NotA);
inv M9_UM9_0_BM18_Xo1(M9_UM9_0_XA3_2, M9_UM9_0_BM18_NotB);
nand2 M9_UM9_0_BM18_Xo2(M9_UM9_0_BM18_NotA, M9_UM9_0_XA3_2, M9_UM9_0_BM18_line2);
nand2 M9_UM9_0_BM18_Xo3(M9_UM9_0_BM18_NotB, M9_UM9_0_XA1_0, M9_UM9_0_BM18_line3);
nand2 M9_UM9_0_BM18_Xo4(M9_UM9_0_BM18_line2, M9_UM9_0_BM18_line3, M9_UM9_0_XA3_0);
inv M9_UM9_0_BM19(M9_UM9_0_XA3_0, M9_temp1bus_2);
inv M9_UM9_0_BM20_Xo0(in270, M9_UM9_0_BM20_NotA);
inv M9_UM9_0_BM20_Xo1(in264, M9_UM9_0_BM20_NotB);
nand2 M9_UM9_0_BM20_Xo2(M9_UM9_0_BM20_NotA, in264, M9_UM9_0_BM20_line2);
nand2 M9_UM9_0_BM20_Xo3(M9_UM9_0_BM20_NotB, in270, M9_UM9_0_BM20_line3);
nand2 M9_UM9_0_BM20_Xo4(M9_UM9_0_BM20_line2, M9_UM9_0_BM20_line3, M9_UM9_0_XB1_0);
inv M9_UM9_0_BM21_Xo0(in257, M9_UM9_0_BM21_NotA);
inv M9_UM9_0_BM21_Xo1(in250, M9_UM9_0_BM21_NotB);
nand2 M9_UM9_0_BM21_Xo2(M9_UM9_0_BM21_NotA, in250, M9_UM9_0_BM21_line2);
nand2 M9_UM9_0_BM21_Xo3(M9_UM9_0_BM21_NotB, in257, M9_UM9_0_BM21_line3);
nand2 M9_UM9_0_BM21_Xo4(M9_UM9_0_BM21_line2, M9_UM9_0_BM21_line3, M9_UM9_0_XB3_2);
inv M9_UM9_0_BM22_Xo0(M9_UM9_0_XB1_0, M9_UM9_0_BM22_NotA);
inv M9_UM9_0_BM22_Xo1(M9_UM9_0_XB3_2, M9_UM9_0_BM22_NotB);
nand2 M9_UM9_0_BM22_Xo2(M9_UM9_0_BM22_NotA, M9_UM9_0_XB3_2, M9_UM9_0_BM22_line2);
nand2 M9_UM9_0_BM22_Xo3(M9_UM9_0_BM22_NotB, M9_UM9_0_XB1_0, M9_UM9_0_BM22_line3);
nand2 M9_UM9_0_BM22_Xo4(M9_UM9_0_BM22_line2, M9_UM9_0_BM22_line3, M9_UM9_0_XB3_0);
inv M9_UM9_0_BM23(M9_UM9_0_XB3_0, M9_temp1bus_3);
nand2 M9_UM9_0_BM24(M9_UM9_0_NotAbus_2, M9_UM9_0_NotAbus_1, M9_UM9_0_NotA1_0);
and2 M9_UM9_0_BM25(in87, M9_UM9_0_NotA1_0, M9_temp2bus_0);
and2 M9_UM9_0_BM26(M9_UM9_0_NotAbus_0, M9_UM9_0_NotA3_1, M9_temp2bus_1);
inv M9_UM9_1(in13, M9_NotCont1);
inv M9_UM9_2(in33, M9_NotCont3);
and3 M9_UM9_3(in1, M9_NotCont1, in20, M9_temp3);
nand2 M9_UM9_4(M9_temp3, in33, M9_ContHi);
nand2 M9_UM9_5(M9_temp3, M9_NotCont3, M9_ContLo);
inv M9_UM9_6_M4b3c_0_Mux3c_0(M9_ContHi, M9_UM9_6_M4b3c_0_NotContHi);
inv M9_UM9_6_M4b3c_0_Mux3c_1(M9_ContLo, M9_UM9_6_M4b3c_0_NotContLo);
and2 M9_UM9_6_M4b3c_0_Mux3c_2(M9_temp1bus_0, M9_UM9_6_M4b3c_0_NotContHi, M9_UM9_6_M4b3c_0_line2);
and2 M9_UM9_6_M4b3c_0_Mux3c_3(M9_temp2bus_0, M9_UM9_6_M4b3c_0_NotContLo, M9_UM9_6_M4b3c_0_line3);
and2 M9_UM9_6_M4b3c_0_Mux3c_4(M9_ContHi, M9_ContLo, M9_UM9_6_M4b3c_0_line4);
and2 M9_UM9_6_M4b3c_0_Mux3c_5(M9_UM9_6_M4b3c_0_line4, in116, M9_UM9_6_M4b3c_0_line5);
or3 M9_UM9_6_M4b3c_0_Mux3c_6(M9_UM9_6_M4b3c_0_line2, M9_UM9_6_M4b3c_0_line3, M9_UM9_6_M4b3c_0_line5, Hbus_0);
inv M9_UM9_6_M4b3c_1_Mux3c_0(M9_ContHi, M9_UM9_6_M4b3c_1_NotContHi);
inv M9_UM9_6_M4b3c_1_Mux3c_1(M9_ContLo, M9_UM9_6_M4b3c_1_NotContLo);
and2 M9_UM9_6_M4b3c_1_Mux3c_2(M9_temp1bus_1, M9_UM9_6_M4b3c_1_NotContHi, M9_UM9_6_M4b3c_1_line2);
and2 M9_UM9_6_M4b3c_1_Mux3c_3(M9_temp2bus_1, M9_UM9_6_M4b3c_1_NotContLo, M9_UM9_6_M4b3c_1_line3);
and2 M9_UM9_6_M4b3c_1_Mux3c_4(M9_ContHi, M9_ContLo, M9_UM9_6_M4b3c_1_line4);
and2 M9_UM9_6_M4b3c_1_Mux3c_5(M9_UM9_6_M4b3c_1_line4, in107, M9_UM9_6_M4b3c_1_line5);
or3 M9_UM9_6_M4b3c_1_Mux3c_6(M9_UM9_6_M4b3c_1_line2, M9_UM9_6_M4b3c_1_line3, M9_UM9_6_M4b3c_1_line5, Hbus_1);
inv M9_UM9_6_M4b3c_2_Mux3c_0(M9_ContHi, M9_UM9_6_M4b3c_2_NotContHi);
inv M9_UM9_6_M4b3c_2_Mux3c_1(M9_ContLo, M9_UM9_6_M4b3c_2_NotContLo);
and2 M9_UM9_6_M4b3c_2_Mux3c_2(M9_temp1bus_2, M9_UM9_6_M4b3c_2_NotContHi, M9_UM9_6_M4b3c_2_line2);
and2 M9_UM9_6_M4b3c_2_Mux3c_3(gnd, M9_UM9_6_M4b3c_2_NotContLo, M9_UM9_6_M4b3c_2_line3);
and2 M9_UM9_6_M4b3c_2_Mux3c_4(M9_ContHi, M9_ContLo, M9_UM9_6_M4b3c_2_line4);
and2 M9_UM9_6_M4b3c_2_Mux3c_5(M9_UM9_6_M4b3c_2_line4, in97, M9_UM9_6_M4b3c_2_line5);
or3 M9_UM9_6_M4b3c_2_Mux3c_6(M9_UM9_6_M4b3c_2_line2, M9_UM9_6_M4b3c_2_line3, M9_UM9_6_M4b3c_2_line5, Hbus_2);
inv M9_UM9_6_M4b3c_3_Mux3c_0(M9_ContHi, M9_UM9_6_M4b3c_3_NotContHi);
inv M9_UM9_6_M4b3c_3_Mux3c_1(M9_ContLo, M9_UM9_6_M4b3c_3_NotContLo);
and2 M9_UM9_6_M4b3c_3_Mux3c_2(M9_temp1bus_3, M9_UM9_6_M4b3c_3_NotContHi, M9_UM9_6_M4b3c_3_line2);
and2 M9_UM9_6_M4b3c_3_Mux3c_3(gnd, M9_UM9_6_M4b3c_3_NotContLo, M9_UM9_6_M4b3c_3_line3);
and2 M9_UM9_6_M4b3c_3_Mux3c_4(M9_ContHi, M9_ContLo, M9_UM9_6_M4b3c_3_line4);
and2 M9_UM9_6_M4b3c_3_Mux3c_5(M9_UM9_6_M4b3c_3_line4, in87, M9_UM9_6_M4b3c_3_line5);
or3 M9_UM9_6_M4b3c_3_Mux3c_6(M9_UM9_6_M4b3c_3_line2, M9_UM9_6_M4b3c_3_line3, M9_UM9_6_M4b3c_3_line5, Hbus_3);
inv M10_UM10_0(in13, M10_NotCont1);
inv M10_UM10_1(in20, M10_NotCont2);
inv M10_UM10_2(in33, M10_NotCont3);
or2 M10_UM10_3(M10_NotCont2, in169, M10_tmp0);
nand3 M10_UM10_4(in1, in13, M10_tmp0, M10_ContHi);
nand3 M10_UM10_5(M10_NotCont1, M10_NotCont2, M10_NotCont3, M10_ContLo1);
nand2 M10_UM10_6(M10_NotCont1, M10_NotCont3, M10_ContLo2);
inv M10_UM10_7_M4b3c_0_Mux3c_0(M10_ContHi, M10_UM10_7_M4b3c_0_NotContHi);
inv M10_UM10_7_M4b3c_0_Mux3c_1(M10_ContLo1, M10_UM10_7_M4b3c_0_NotContLo);
and2 M10_UM10_7_M4b3c_0_Mux3c_2(Shiftbus_0, M10_UM10_7_M4b3c_0_NotContHi, M10_UM10_7_M4b3c_0_line2);
and2 M10_UM10_7_M4b3c_0_Mux3c_3(XPbus_0, M10_UM10_7_M4b3c_0_NotContLo, M10_UM10_7_M4b3c_0_line3);
and2 M10_UM10_7_M4b3c_0_Mux3c_4(M10_ContHi, M10_ContLo1, M10_UM10_7_M4b3c_0_line4);
and2 M10_UM10_7_M4b3c_0_Mux3c_5(M10_UM10_7_M4b3c_0_line4, Hbus_0, M10_UM10_7_M4b3c_0_line5);
or3 M10_UM10_7_M4b3c_0_Mux3c_6(M10_UM10_7_M4b3c_0_line2, M10_UM10_7_M4b3c_0_line3, M10_UM10_7_M4b3c_0_line5, Wbus_0);
inv M10_UM10_7_M4b3c_1_Mux3c_0(M10_ContHi, M10_UM10_7_M4b3c_1_NotContHi);
inv M10_UM10_7_M4b3c_1_Mux3c_1(M10_ContLo1, M10_UM10_7_M4b3c_1_NotContLo);
and2 M10_UM10_7_M4b3c_1_Mux3c_2(Shiftbus_1, M10_UM10_7_M4b3c_1_NotContHi, M10_UM10_7_M4b3c_1_line2);
and2 M10_UM10_7_M4b3c_1_Mux3c_3(XPbus_1, M10_UM10_7_M4b3c_1_NotContLo, M10_UM10_7_M4b3c_1_line3);
and2 M10_UM10_7_M4b3c_1_Mux3c_4(M10_ContHi, M10_ContLo1, M10_UM10_7_M4b3c_1_line4);
and2 M10_UM10_7_M4b3c_1_Mux3c_5(M10_UM10_7_M4b3c_1_line4, Hbus_1, M10_UM10_7_M4b3c_1_line5);
or3 M10_UM10_7_M4b3c_1_Mux3c_6(M10_UM10_7_M4b3c_1_line2, M10_UM10_7_M4b3c_1_line3, M10_UM10_7_M4b3c_1_line5, Wbus_1);
inv M10_UM10_7_M4b3c_2_Mux3c_0(M10_ContHi, M10_UM10_7_M4b3c_2_NotContHi);
inv M10_UM10_7_M4b3c_2_Mux3c_1(M10_ContLo1, M10_UM10_7_M4b3c_2_NotContLo);
and2 M10_UM10_7_M4b3c_2_Mux3c_2(Shiftbus_2, M10_UM10_7_M4b3c_2_NotContHi, M10_UM10_7_M4b3c_2_line2);
and2 M10_UM10_7_M4b3c_2_Mux3c_3(XPbus_2, M10_UM10_7_M4b3c_2_NotContLo, M10_UM10_7_M4b3c_2_line3);
and2 M10_UM10_7_M4b3c_2_Mux3c_4(M10_ContHi, M10_ContLo1, M10_UM10_7_M4b3c_2_line4);
and2 M10_UM10_7_M4b3c_2_Mux3c_5(M10_UM10_7_M4b3c_2_line4, Hbus_2, M10_UM10_7_M4b3c_2_line5);
or3 M10_UM10_7_M4b3c_2_Mux3c_6(M10_UM10_7_M4b3c_2_line2, M10_UM10_7_M4b3c_2_line3, M10_UM10_7_M4b3c_2_line5, Wbus_2);
inv M10_UM10_7_M4b3c_3_Mux3c_0(M10_ContHi, M10_UM10_7_M4b3c_3_NotContHi);
inv M10_UM10_7_M4b3c_3_Mux3c_1(M10_ContLo1, M10_UM10_7_M4b3c_3_NotContLo);
and2 M10_UM10_7_M4b3c_3_Mux3c_2(Shiftbus_3, M10_UM10_7_M4b3c_3_NotContHi, M10_UM10_7_M4b3c_3_line2);
and2 M10_UM10_7_M4b3c_3_Mux3c_3(XPbus_3, M10_UM10_7_M4b3c_3_NotContLo, M10_UM10_7_M4b3c_3_line3);
and2 M10_UM10_7_M4b3c_3_Mux3c_4(M10_ContHi, M10_ContLo1, M10_UM10_7_M4b3c_3_line4);
and2 M10_UM10_7_M4b3c_3_Mux3c_5(M10_UM10_7_M4b3c_3_line4, Hbus_3, M10_UM10_7_M4b3c_3_line5);
or3 M10_UM10_7_M4b3c_3_Mux3c_6(M10_UM10_7_M4b3c_3_line2, M10_UM10_7_M4b3c_3_line3, M10_UM10_7_M4b3c_3_line5, Wbus_3);
inv M10_UM10_8_M4b3c_0_Mux3c_0(M10_ContHi, M10_UM10_8_M4b3c_0_NotContHi);
inv M10_UM10_8_M4b3c_0_Mux3c_1(M10_ContLo2, M10_UM10_8_M4b3c_0_NotContLo);
and2 M10_UM10_8_M4b3c_0_Mux3c_2(Shiftbus_4, M10_UM10_8_M4b3c_0_NotContHi, M10_UM10_8_M4b3c_0_line2);
and2 M10_UM10_8_M4b3c_0_Mux3c_3(XPbus_4, M10_UM10_8_M4b3c_0_NotContLo, M10_UM10_8_M4b3c_0_line3);
and2 M10_UM10_8_M4b3c_0_Mux3c_4(M10_ContHi, M10_ContLo2, M10_UM10_8_M4b3c_0_line4);
and2 M10_UM10_8_M4b3c_0_Mux3c_5(M10_UM10_8_M4b3c_0_line4, in77, M10_UM10_8_M4b3c_0_line5);
or3 M10_UM10_8_M4b3c_0_Mux3c_6(M10_UM10_8_M4b3c_0_line2, M10_UM10_8_M4b3c_0_line3, M10_UM10_8_M4b3c_0_line5, Wbus_4);
inv M10_UM10_8_M4b3c_1_Mux3c_0(M10_ContHi, M10_UM10_8_M4b3c_1_NotContHi);
inv M10_UM10_8_M4b3c_1_Mux3c_1(M10_ContLo2, M10_UM10_8_M4b3c_1_NotContLo);
and2 M10_UM10_8_M4b3c_1_Mux3c_2(Shiftbus_5, M10_UM10_8_M4b3c_1_NotContHi, M10_UM10_8_M4b3c_1_line2);
and2 M10_UM10_8_M4b3c_1_Mux3c_3(XPbus_5, M10_UM10_8_M4b3c_1_NotContLo, M10_UM10_8_M4b3c_1_line3);
and2 M10_UM10_8_M4b3c_1_Mux3c_4(M10_ContHi, M10_ContLo2, M10_UM10_8_M4b3c_1_line4);
and2 M10_UM10_8_M4b3c_1_Mux3c_5(M10_UM10_8_M4b3c_1_line4, in68, M10_UM10_8_M4b3c_1_line5);
or3 M10_UM10_8_M4b3c_1_Mux3c_6(M10_UM10_8_M4b3c_1_line2, M10_UM10_8_M4b3c_1_line3, M10_UM10_8_M4b3c_1_line5, Wbus_5);
inv M10_UM10_8_M4b3c_2_Mux3c_0(M10_ContHi, M10_UM10_8_M4b3c_2_NotContHi);
inv M10_UM10_8_M4b3c_2_Mux3c_1(M10_ContLo2, M10_UM10_8_M4b3c_2_NotContLo);
and2 M10_UM10_8_M4b3c_2_Mux3c_2(Shiftbus_6, M10_UM10_8_M4b3c_2_NotContHi, M10_UM10_8_M4b3c_2_line2);
and2 M10_UM10_8_M4b3c_2_Mux3c_3(XPbus_6, M10_UM10_8_M4b3c_2_NotContLo, M10_UM10_8_M4b3c_2_line3);
and2 M10_UM10_8_M4b3c_2_Mux3c_4(M10_ContHi, M10_ContLo2, M10_UM10_8_M4b3c_2_line4);
and2 M10_UM10_8_M4b3c_2_Mux3c_5(M10_UM10_8_M4b3c_2_line4, in58, M10_UM10_8_M4b3c_2_line5);
or3 M10_UM10_8_M4b3c_2_Mux3c_6(M10_UM10_8_M4b3c_2_line2, M10_UM10_8_M4b3c_2_line3, M10_UM10_8_M4b3c_2_line5, Wbus_6);
inv M10_UM10_8_M4b3c_3_Mux3c_0(M10_ContHi, M10_UM10_8_M4b3c_3_NotContHi);
inv M10_UM10_8_M4b3c_3_Mux3c_1(M10_ContLo2, M10_UM10_8_M4b3c_3_NotContLo);
and2 M10_UM10_8_M4b3c_3_Mux3c_2(Shiftbus_7, M10_UM10_8_M4b3c_3_NotContHi, M10_UM10_8_M4b3c_3_line2);
and2 M10_UM10_8_M4b3c_3_Mux3c_3(XPbus_7, M10_UM10_8_M4b3c_3_NotContLo, M10_UM10_8_M4b3c_3_line3);
and2 M10_UM10_8_M4b3c_3_Mux3c_4(M10_ContHi, M10_ContLo2, M10_UM10_8_M4b3c_3_line4);
and2 M10_UM10_8_M4b3c_3_Mux3c_5(M10_UM10_8_M4b3c_3_line4, in50, M10_UM10_8_M4b3c_3_line5);
or3 M10_UM10_8_M4b3c_3_Mux3c_6(M10_UM10_8_M4b3c_3_line2, M10_UM10_8_M4b3c_3_line3, M10_UM10_8_M4b3c_3_line5, Wbus_7);
inv M11_UM11_0(in13, M11_NotCont1);
inv M11_UM11_1(in20, M11_NotCont2);
inv M11_UM11_2(in41, M11_NotCont5);
nand3 M11_UM11_3(in13, M11_NotCont2, in45, M11_tmp0);
and2 M11_UM11_4(in1, M11_tmp0, M11_ContHi);
nand4 M11_UM11_5(in1, M11_NotCont1, in20, M11_NotCont5, M11_ContLo);
inv M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_0_M4b3c_0_NotContHi);
inv M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_0_NotContLo);
and2 M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_2(Funcbus_0, M11_UM11_7_M8b3c_0_M4b3c_0_NotContHi, M11_UM11_7_M8b3c_0_M4b3c_0_line2);
and2 M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_3(Funcbus_0, M11_UM11_7_M8b3c_0_M4b3c_0_NotContLo, M11_UM11_7_M8b3c_0_M4b3c_0_line3);
and2 M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_0_line4);
and2 M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_5(M11_UM11_7_M8b3c_0_M4b3c_0_line4, Wbus_0, M11_UM11_7_M8b3c_0_M4b3c_0_line5);
or3 M11_UM11_7_M8b3c_0_M4b3c_0_Mux3c_6(M11_UM11_7_M8b3c_0_M4b3c_0_line2, M11_UM11_7_M8b3c_0_M4b3c_0_line3, M11_UM11_7_M8b3c_0_M4b3c_0_line5, out396);
inv M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_0_M4b3c_1_NotContHi);
inv M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_1_NotContLo);
and2 M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_2(Funcbus_1, M11_UM11_7_M8b3c_0_M4b3c_1_NotContHi, M11_UM11_7_M8b3c_0_M4b3c_1_line2);
and2 M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_3(F_BCDbus_1, M11_UM11_7_M8b3c_0_M4b3c_1_NotContLo, M11_UM11_7_M8b3c_0_M4b3c_1_line3);
and2 M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_1_line4);
and2 M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_5(M11_UM11_7_M8b3c_0_M4b3c_1_line4, Wbus_1, M11_UM11_7_M8b3c_0_M4b3c_1_line5);
or3 M11_UM11_7_M8b3c_0_M4b3c_1_Mux3c_6(M11_UM11_7_M8b3c_0_M4b3c_1_line2, M11_UM11_7_M8b3c_0_M4b3c_1_line3, M11_UM11_7_M8b3c_0_M4b3c_1_line5, out393);
inv M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_0_M4b3c_2_NotContHi);
inv M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_2_NotContLo);
and2 M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_2(Funcbus_2, M11_UM11_7_M8b3c_0_M4b3c_2_NotContHi, M11_UM11_7_M8b3c_0_M4b3c_2_line2);
and2 M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_3(F_BCDbus_2, M11_UM11_7_M8b3c_0_M4b3c_2_NotContLo, M11_UM11_7_M8b3c_0_M4b3c_2_line3);
and2 M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_2_line4);
and2 M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_5(M11_UM11_7_M8b3c_0_M4b3c_2_line4, Wbus_2, M11_UM11_7_M8b3c_0_M4b3c_2_line5);
or3 M11_UM11_7_M8b3c_0_M4b3c_2_Mux3c_6(M11_UM11_7_M8b3c_0_M4b3c_2_line2, M11_UM11_7_M8b3c_0_M4b3c_2_line3, M11_UM11_7_M8b3c_0_M4b3c_2_line5, out390);
inv M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_0_M4b3c_3_NotContHi);
inv M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_3_NotContLo);
and2 M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_2(Funcbus_3, M11_UM11_7_M8b3c_0_M4b3c_3_NotContHi, M11_UM11_7_M8b3c_0_M4b3c_3_line2);
and2 M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_3(F_BCDbus_3, M11_UM11_7_M8b3c_0_M4b3c_3_NotContLo, M11_UM11_7_M8b3c_0_M4b3c_3_line3);
and2 M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_0_M4b3c_3_line4);
and2 M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_5(M11_UM11_7_M8b3c_0_M4b3c_3_line4, Wbus_3, M11_UM11_7_M8b3c_0_M4b3c_3_line5);
or3 M11_UM11_7_M8b3c_0_M4b3c_3_Mux3c_6(M11_UM11_7_M8b3c_0_M4b3c_3_line2, M11_UM11_7_M8b3c_0_M4b3c_3_line3, M11_UM11_7_M8b3c_0_M4b3c_3_line5, out387);
inv M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_1_M4b3c_0_NotContHi);
inv M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_0_NotContLo);
and2 M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_2(Funcbus_4, M11_UM11_7_M8b3c_1_M4b3c_0_NotContHi, M11_UM11_7_M8b3c_1_M4b3c_0_line2);
and2 M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_3(Funcbus_4, M11_UM11_7_M8b3c_1_M4b3c_0_NotContLo, M11_UM11_7_M8b3c_1_M4b3c_0_line3);
and2 M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_0_line4);
and2 M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_5(M11_UM11_7_M8b3c_1_M4b3c_0_line4, Wbus_4, M11_UM11_7_M8b3c_1_M4b3c_0_line5);
or3 M11_UM11_7_M8b3c_1_M4b3c_0_Mux3c_6(M11_UM11_7_M8b3c_1_M4b3c_0_line2, M11_UM11_7_M8b3c_1_M4b3c_0_line3, M11_UM11_7_M8b3c_1_M4b3c_0_line5, out384);
inv M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_1_M4b3c_1_NotContHi);
inv M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_1_NotContLo);
and2 M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_2(Funcbus_5, M11_UM11_7_M8b3c_1_M4b3c_1_NotContHi, M11_UM11_7_M8b3c_1_M4b3c_1_line2);
and2 M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_3(F_BCDbus_5, M11_UM11_7_M8b3c_1_M4b3c_1_NotContLo, M11_UM11_7_M8b3c_1_M4b3c_1_line3);
and2 M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_1_line4);
and2 M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_5(M11_UM11_7_M8b3c_1_M4b3c_1_line4, Wbus_5, M11_UM11_7_M8b3c_1_M4b3c_1_line5);
or3 M11_UM11_7_M8b3c_1_M4b3c_1_Mux3c_6(M11_UM11_7_M8b3c_1_M4b3c_1_line2, M11_UM11_7_M8b3c_1_M4b3c_1_line3, M11_UM11_7_M8b3c_1_M4b3c_1_line5, out381);
inv M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_1_M4b3c_2_NotContHi);
inv M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_2_NotContLo);
and2 M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_2(Funcbus_6, M11_UM11_7_M8b3c_1_M4b3c_2_NotContHi, M11_UM11_7_M8b3c_1_M4b3c_2_line2);
and2 M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_3(F_BCDbus_6, M11_UM11_7_M8b3c_1_M4b3c_2_NotContLo, M11_UM11_7_M8b3c_1_M4b3c_2_line3);
and2 M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_2_line4);
and2 M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_5(M11_UM11_7_M8b3c_1_M4b3c_2_line4, Wbus_6, M11_UM11_7_M8b3c_1_M4b3c_2_line5);
or3 M11_UM11_7_M8b3c_1_M4b3c_2_Mux3c_6(M11_UM11_7_M8b3c_1_M4b3c_2_line2, M11_UM11_7_M8b3c_1_M4b3c_2_line3, M11_UM11_7_M8b3c_1_M4b3c_2_line5, out378);
inv M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_0(M11_ContHi, M11_UM11_7_M8b3c_1_M4b3c_3_NotContHi);
inv M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_1(M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_3_NotContLo);
and2 M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_2(Funcbus_7, M11_UM11_7_M8b3c_1_M4b3c_3_NotContHi, M11_UM11_7_M8b3c_1_M4b3c_3_line2);
and2 M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_3(F_BCDbus_7, M11_UM11_7_M8b3c_1_M4b3c_3_NotContLo, M11_UM11_7_M8b3c_1_M4b3c_3_line3);
and2 M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_4(M11_ContHi, M11_ContLo, M11_UM11_7_M8b3c_1_M4b3c_3_line4);
and2 M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_5(M11_UM11_7_M8b3c_1_M4b3c_3_line4, Wbus_7, M11_UM11_7_M8b3c_1_M4b3c_3_line5);
or3 M11_UM11_7_M8b3c_1_M4b3c_3_Mux3c_6(M11_UM11_7_M8b3c_1_M4b3c_3_line2, M11_UM11_7_M8b3c_1_M4b3c_3_line3, M11_UM11_7_M8b3c_1_M4b3c_3_line5, out375);
inv M12_UM12_0_Inv8_0_Inv4_0(out396, M12_Not_Zbus_0);
inv M12_UM12_0_Inv8_0_Inv4_1(out393, M12_Not_Zbus_1);
inv M12_UM12_0_Inv8_0_Inv4_2(out390, M12_Not_Zbus_2);
inv M12_UM12_0_Inv8_0_Inv4_3(out387, M12_Not_Zbus_3);
inv M12_UM12_0_Inv8_1_Inv4_0(out384, M12_Not_Zbus_4);
inv M12_UM12_0_Inv8_1_Inv4_1(out381, M12_Not_Zbus_5);
inv M12_UM12_0_Inv8_1_Inv4_2(out378, M12_Not_Zbus_6);
inv M12_UM12_0_Inv8_1_Inv4_3(out375, M12_Not_Zbus_7);
and4 M12_UM12_1(M12_Not_Zbus_0, M12_Not_Zbus_1, M12_Not_Zbus_2, M12_Not_Zbus_3, M12_ZeroZ_Lo);
and4 M12_UM12_2(M12_Not_Zbus_4, M12_Not_Zbus_5, M12_Not_Zbus_6, M12_Not_Zbus_7, M12_ZeroZ_Hi);
and2 M12_UM12_3(M12_ZeroZ_Lo, M12_ZeroZ_Hi, M12_ZeroZ);
inv M12_UM12_4(M12_ZeroZ, out407);
inv M12_UM12_5(in213, M12_NotCont8);
or2 M12_UM12_6(M12_NotCont8, in343, M12_ContFlag);
inv M12_UM12_7(M12_ContFlag, M12_NotContFlag);
and3 M12_UM12_8(M12_Not_Zbus_6, M12_Not_Zbus_7, M12_NotContFlag, M12_tmp0);
nor2 M12_UM12_9(M12_tmp0, M12_ZeroZ, M12_tmp1);
nand2 M12_UM12_10(in213, M12_tmp1, out409);
inv M12_UM12_11_PT1_Xo0(in116, M12_UM12_11_PT1_NotA);
inv M12_UM12_11_PT1_Xo1(in107, M12_UM12_11_PT1_NotB);
nand2 M12_UM12_11_PT1_Xo2(M12_UM12_11_PT1_NotA, in107, M12_UM12_11_PT1_line2);
nand2 M12_UM12_11_PT1_Xo3(M12_UM12_11_PT1_NotB, in116, M12_UM12_11_PT1_line3);
nand2 M12_UM12_11_PT1_Xo4(M12_UM12_11_PT1_line2, M12_UM12_11_PT1_line3, M12_UM12_11_line1);
inv M12_UM12_11_PT2_Xo0(in97, M12_UM12_11_PT2_NotA);
inv M12_UM12_11_PT2_Xo1(in87, M12_UM12_11_PT2_NotB);
nand2 M12_UM12_11_PT2_Xo2(M12_UM12_11_PT2_NotA, in87, M12_UM12_11_PT2_line2);
nand2 M12_UM12_11_PT2_Xo3(M12_UM12_11_PT2_NotB, in97, M12_UM12_11_PT2_line3);
nand2 M12_UM12_11_PT2_Xo4(M12_UM12_11_PT2_line2, M12_UM12_11_PT2_line3, M12_UM12_11_line2);
inv M12_UM12_11_PT3_Xo0(in77, M12_UM12_11_PT3_NotA);
inv M12_UM12_11_PT3_Xo1(in68, M12_UM12_11_PT3_NotB);
nand2 M12_UM12_11_PT3_Xo2(M12_UM12_11_PT3_NotA, in68, M12_UM12_11_PT3_line2);
nand2 M12_UM12_11_PT3_Xo3(M12_UM12_11_PT3_NotB, in77, M12_UM12_11_PT3_line3);
nand2 M12_UM12_11_PT3_Xo4(M12_UM12_11_PT3_line2, M12_UM12_11_PT3_line3, M12_UM12_11_line3);
inv M12_UM12_11_PT4_Xo0(in58, M12_UM12_11_PT4_NotA);
inv M12_UM12_11_PT4_Xo1(in50, M12_UM12_11_PT4_NotB);
nand2 M12_UM12_11_PT4_Xo2(M12_UM12_11_PT4_NotA, in50, M12_UM12_11_PT4_line2);
nand2 M12_UM12_11_PT4_Xo3(M12_UM12_11_PT4_NotB, in58, M12_UM12_11_PT4_line3);
nand2 M12_UM12_11_PT4_Xo4(M12_UM12_11_PT4_line2, M12_UM12_11_PT4_line3, M12_UM12_11_line4);
inv M12_UM12_11_PT5_Xo0(M12_UM12_11_line1, M12_UM12_11_PT5_NotA);
inv M12_UM12_11_PT5_Xo1(M12_UM12_11_line2, M12_UM12_11_PT5_NotB);
nand2 M12_UM12_11_PT5_Xo2(M12_UM12_11_PT5_NotA, M12_UM12_11_line2, M12_UM12_11_PT5_line2);
nand2 M12_UM12_11_PT5_Xo3(M12_UM12_11_PT5_NotB, M12_UM12_11_line1, M12_UM12_11_PT5_line3);
nand2 M12_UM12_11_PT5_Xo4(M12_UM12_11_PT5_line2, M12_UM12_11_PT5_line3, M12_UM12_11_line5);
inv M12_UM12_11_PT6_Xo0(M12_UM12_11_line3, M12_UM12_11_PT6_NotA);
inv M12_UM12_11_PT6_Xo1(M12_UM12_11_line4, M12_UM12_11_PT6_NotB);
nand2 M12_UM12_11_PT6_Xo2(M12_UM12_11_PT6_NotA, M12_UM12_11_line4, M12_UM12_11_PT6_line2);
nand2 M12_UM12_11_PT6_Xo3(M12_UM12_11_PT6_NotB, M12_UM12_11_line3, M12_UM12_11_PT6_line3);
nand2 M12_UM12_11_PT6_Xo4(M12_UM12_11_PT6_line2, M12_UM12_11_PT6_line3, M12_UM12_11_line6);
inv M12_UM12_11_PT7_Xo0(M12_UM12_11_line5, M12_UM12_11_PT7_NotA);
inv M12_UM12_11_PT7_Xo1(M12_UM12_11_line6, M12_UM12_11_PT7_NotB);
nand2 M12_UM12_11_PT7_Xo2(M12_UM12_11_PT7_NotA, M12_UM12_11_line6, M12_UM12_11_PT7_line2);
nand2 M12_UM12_11_PT7_Xo3(M12_UM12_11_PT7_NotB, M12_UM12_11_line5, M12_UM12_11_PT7_line3);
nand2 M12_UM12_11_PT7_Xo4(M12_UM12_11_PT7_line2, M12_UM12_11_PT7_line3, M12_EvenParA);
inv M12_UM12_12_PT1_Xo0(in270, M12_UM12_12_PT1_NotA);
inv M12_UM12_12_PT1_Xo1(in264, M12_UM12_12_PT1_NotB);
nand2 M12_UM12_12_PT1_Xo2(M12_UM12_12_PT1_NotA, in264, M12_UM12_12_PT1_line2);
nand2 M12_UM12_12_PT1_Xo3(M12_UM12_12_PT1_NotB, in270, M12_UM12_12_PT1_line3);
nand2 M12_UM12_12_PT1_Xo4(M12_UM12_12_PT1_line2, M12_UM12_12_PT1_line3, M12_UM12_12_line1);
inv M12_UM12_12_PT2_Xo0(in257, M12_UM12_12_PT2_NotA);
inv M12_UM12_12_PT2_Xo1(in250, M12_UM12_12_PT2_NotB);
nand2 M12_UM12_12_PT2_Xo2(M12_UM12_12_PT2_NotA, in250, M12_UM12_12_PT2_line2);
nand2 M12_UM12_12_PT2_Xo3(M12_UM12_12_PT2_NotB, in257, M12_UM12_12_PT2_line3);
nand2 M12_UM12_12_PT2_Xo4(M12_UM12_12_PT2_line2, M12_UM12_12_PT2_line3, M12_UM12_12_line2);
inv M12_UM12_12_PT3_Xo0(in244, M12_UM12_12_PT3_NotA);
inv M12_UM12_12_PT3_Xo1(in238, M12_UM12_12_PT3_NotB);
nand2 M12_UM12_12_PT3_Xo2(M12_UM12_12_PT3_NotA, in238, M12_UM12_12_PT3_line2);
nand2 M12_UM12_12_PT3_Xo3(M12_UM12_12_PT3_NotB, in244, M12_UM12_12_PT3_line3);
nand2 M12_UM12_12_PT3_Xo4(M12_UM12_12_PT3_line2, M12_UM12_12_PT3_line3, M12_UM12_12_line3);
inv M12_UM12_12_PT4_Xo0(in232, M12_UM12_12_PT4_NotA);
inv M12_UM12_12_PT4_Xo1(in226, M12_UM12_12_PT4_NotB);
nand2 M12_UM12_12_PT4_Xo2(M12_UM12_12_PT4_NotA, in226, M12_UM12_12_PT4_line2);
nand2 M12_UM12_12_PT4_Xo3(M12_UM12_12_PT4_NotB, in232, M12_UM12_12_PT4_line3);
nand2 M12_UM12_12_PT4_Xo4(M12_UM12_12_PT4_line2, M12_UM12_12_PT4_line3, M12_UM12_12_line4);
inv M12_UM12_12_PT5_Xo0(M12_UM12_12_line1, M12_UM12_12_PT5_NotA);
inv M12_UM12_12_PT5_Xo1(M12_UM12_12_line2, M12_UM12_12_PT5_NotB);
nand2 M12_UM12_12_PT5_Xo2(M12_UM12_12_PT5_NotA, M12_UM12_12_line2, M12_UM12_12_PT5_line2);
nand2 M12_UM12_12_PT5_Xo3(M12_UM12_12_PT5_NotB, M12_UM12_12_line1, M12_UM12_12_PT5_line3);
nand2 M12_UM12_12_PT5_Xo4(M12_UM12_12_PT5_line2, M12_UM12_12_PT5_line3, M12_UM12_12_line5);
inv M12_UM12_12_PT6_Xo0(M12_UM12_12_line3, M12_UM12_12_PT6_NotA);
inv M12_UM12_12_PT6_Xo1(M12_UM12_12_line4, M12_UM12_12_PT6_NotB);
nand2 M12_UM12_12_PT6_Xo2(M12_UM12_12_PT6_NotA, M12_UM12_12_line4, M12_UM12_12_PT6_line2);
nand2 M12_UM12_12_PT6_Xo3(M12_UM12_12_PT6_NotB, M12_UM12_12_line3, M12_UM12_12_PT6_line3);
nand2 M12_UM12_12_PT6_Xo4(M12_UM12_12_PT6_line2, M12_UM12_12_PT6_line3, M12_UM12_12_line6);
inv M12_UM12_12_PT7_Xo0(M12_UM12_12_line5, M12_UM12_12_PT7_NotA);
inv M12_UM12_12_PT7_Xo1(M12_UM12_12_line6, M12_UM12_12_PT7_NotB);
nand2 M12_UM12_12_PT7_Xo2(M12_UM12_12_PT7_NotA, M12_UM12_12_line6, M12_UM12_12_PT7_line2);
nand2 M12_UM12_12_PT7_Xo3(M12_UM12_12_PT7_NotB, M12_UM12_12_line5, M12_UM12_12_PT7_line3);
nand2 M12_UM12_12_PT7_Xo4(M12_UM12_12_PT7_line2, M12_UM12_12_PT7_line3, M12_EvenParB);
inv M12_UM12_13_PT1_Xo0(out396, M12_UM12_13_PT1_NotA);
inv M12_UM12_13_PT1_Xo1(out393, M12_UM12_13_PT1_NotB);
nand2 M12_UM12_13_PT1_Xo2(M12_UM12_13_PT1_NotA, out393, M12_UM12_13_PT1_line2);
nand2 M12_UM12_13_PT1_Xo3(M12_UM12_13_PT1_NotB, out396, M12_UM12_13_PT1_line3);
nand2 M12_UM12_13_PT1_Xo4(M12_UM12_13_PT1_line2, M12_UM12_13_PT1_line3, M12_UM12_13_line1);
inv M12_UM12_13_PT2_Xo0(out390, M12_UM12_13_PT2_NotA);
inv M12_UM12_13_PT2_Xo1(out387, M12_UM12_13_PT2_NotB);
nand2 M12_UM12_13_PT2_Xo2(M12_UM12_13_PT2_NotA, out387, M12_UM12_13_PT2_line2);
nand2 M12_UM12_13_PT2_Xo3(M12_UM12_13_PT2_NotB, out390, M12_UM12_13_PT2_line3);
nand2 M12_UM12_13_PT2_Xo4(M12_UM12_13_PT2_line2, M12_UM12_13_PT2_line3, M12_UM12_13_line2);
inv M12_UM12_13_PT3_Xo0(out384, M12_UM12_13_PT3_NotA);
inv M12_UM12_13_PT3_Xo1(out381, M12_UM12_13_PT3_NotB);
nand2 M12_UM12_13_PT3_Xo2(M12_UM12_13_PT3_NotA, out381, M12_UM12_13_PT3_line2);
nand2 M12_UM12_13_PT3_Xo3(M12_UM12_13_PT3_NotB, out384, M12_UM12_13_PT3_line3);
nand2 M12_UM12_13_PT3_Xo4(M12_UM12_13_PT3_line2, M12_UM12_13_PT3_line3, M12_UM12_13_line3);
inv M12_UM12_13_PT4_Xo0(out378, M12_UM12_13_PT4_NotA);
inv M12_UM12_13_PT4_Xo1(out375, M12_UM12_13_PT4_NotB);
nand2 M12_UM12_13_PT4_Xo2(M12_UM12_13_PT4_NotA, out375, M12_UM12_13_PT4_line2);
nand2 M12_UM12_13_PT4_Xo3(M12_UM12_13_PT4_NotB, out378, M12_UM12_13_PT4_line3);
nand2 M12_UM12_13_PT4_Xo4(M12_UM12_13_PT4_line2, M12_UM12_13_PT4_line3, M12_UM12_13_line4);
inv M12_UM12_13_PT5_Xo0(M12_UM12_13_line1, M12_UM12_13_PT5_NotA);
inv M12_UM12_13_PT5_Xo1(M12_UM12_13_line2, M12_UM12_13_PT5_NotB);
nand2 M12_UM12_13_PT5_Xo2(M12_UM12_13_PT5_NotA, M12_UM12_13_line2, M12_UM12_13_PT5_line2);
nand2 M12_UM12_13_PT5_Xo3(M12_UM12_13_PT5_NotB, M12_UM12_13_line1, M12_UM12_13_PT5_line3);
nand2 M12_UM12_13_PT5_Xo4(M12_UM12_13_PT5_line2, M12_UM12_13_PT5_line3, M12_UM12_13_line5);
inv M12_UM12_13_PT6_Xo0(M12_UM12_13_line3, M12_UM12_13_PT6_NotA);
inv M12_UM12_13_PT6_Xo1(M12_UM12_13_line4, M12_UM12_13_PT6_NotB);
nand2 M12_UM12_13_PT6_Xo2(M12_UM12_13_PT6_NotA, M12_UM12_13_line4, M12_UM12_13_PT6_line2);
nand2 M12_UM12_13_PT6_Xo3(M12_UM12_13_PT6_NotB, M12_UM12_13_line3, M12_UM12_13_PT6_line3);
nand2 M12_UM12_13_PT6_Xo4(M12_UM12_13_PT6_line2, M12_UM12_13_PT6_line3, M12_UM12_13_line6);
inv M12_UM12_13_PT7_Xo0(M12_UM12_13_line5, M12_UM12_13_PT7_NotA);
inv M12_UM12_13_PT7_Xo1(M12_UM12_13_line6, M12_UM12_13_PT7_NotB);
nand2 M12_UM12_13_PT7_Xo2(M12_UM12_13_PT7_NotA, M12_UM12_13_line6, M12_UM12_13_PT7_line2);
nand2 M12_UM12_13_PT7_Xo3(M12_UM12_13_PT7_NotB, M12_UM12_13_line5, M12_UM12_13_PT7_line3);
nand2 M12_UM12_13_PT7_Xo4(M12_UM12_13_PT7_line2, M12_UM12_13_PT7_line3, M12_EvenParZ);
and2 M12_UM12_14(M12_NotContFlag, in2897, M12_ContPar);
and2 M12_UM12_15(M12_ContFlag, out375, M12_PZ7);
and2 M12_UM12_16(M12_ContFlag, out378, M12_PZ6);
inv M12_UM12_17_PT1_Xo0(out396, M12_UM12_17_PT1_NotA);
inv M12_UM12_17_PT1_Xo1(out393, M12_UM12_17_PT1_NotB);
nand2 M12_UM12_17_PT1_Xo2(M12_UM12_17_PT1_NotA, out393, M12_UM12_17_PT1_line2);
nand2 M12_UM12_17_PT1_Xo3(M12_UM12_17_PT1_NotB, out396, M12_UM12_17_PT1_line3);
nand2 M12_UM12_17_PT1_Xo4(M12_UM12_17_PT1_line2, M12_UM12_17_PT1_line3, M12_UM12_17_line1);
inv M12_UM12_17_PT2_Xo0(out390, M12_UM12_17_PT2_NotA);
inv M12_UM12_17_PT2_Xo1(out387, M12_UM12_17_PT2_NotB);
nand2 M12_UM12_17_PT2_Xo2(M12_UM12_17_PT2_NotA, out387, M12_UM12_17_PT2_line2);
nand2 M12_UM12_17_PT2_Xo3(M12_UM12_17_PT2_NotB, out390, M12_UM12_17_PT2_line3);
nand2 M12_UM12_17_PT2_Xo4(M12_UM12_17_PT2_line2, M12_UM12_17_PT2_line3, M12_UM12_17_line2);
inv M12_UM12_17_PT3_Xo0(out384, M12_UM12_17_PT3_NotA);
inv M12_UM12_17_PT3_Xo1(out381, M12_UM12_17_PT3_NotB);
nand2 M12_UM12_17_PT3_Xo2(M12_UM12_17_PT3_NotA, out381, M12_UM12_17_PT3_line2);
nand2 M12_UM12_17_PT3_Xo3(M12_UM12_17_PT3_NotB, out384, M12_UM12_17_PT3_line3);
nand2 M12_UM12_17_PT3_Xo4(M12_UM12_17_PT3_line2, M12_UM12_17_PT3_line3, M12_UM12_17_line3);
inv M12_UM12_17_PT4_Xo0(M12_PZ6, M12_UM12_17_PT4_NotA);
inv M12_UM12_17_PT4_Xo1(M12_PZ7, M12_UM12_17_PT4_NotB);
nand2 M12_UM12_17_PT4_Xo2(M12_UM12_17_PT4_NotA, M12_PZ7, M12_UM12_17_PT4_line2);
nand2 M12_UM12_17_PT4_Xo3(M12_UM12_17_PT4_NotB, M12_PZ6, M12_UM12_17_PT4_line3);
nand2 M12_UM12_17_PT4_Xo4(M12_UM12_17_PT4_line2, M12_UM12_17_PT4_line3, M12_UM12_17_line4);
inv M12_UM12_17_PT5_Xo0(M12_UM12_17_line1, M12_UM12_17_PT5_NotA);
inv M12_UM12_17_PT5_Xo1(M12_UM12_17_line2, M12_UM12_17_PT5_NotB);
nand2 M12_UM12_17_PT5_Xo2(M12_UM12_17_PT5_NotA, M12_UM12_17_line2, M12_UM12_17_PT5_line2);
nand2 M12_UM12_17_PT5_Xo3(M12_UM12_17_PT5_NotB, M12_UM12_17_line1, M12_UM12_17_PT5_line3);
nand2 M12_UM12_17_PT5_Xo4(M12_UM12_17_PT5_line2, M12_UM12_17_PT5_line3, M12_UM12_17_line5);
inv M12_UM12_17_PT6_Xo3_0(M12_UM12_17_line3, M12_UM12_17_PT6_NotA);
inv M12_UM12_17_PT6_Xo3_1(M12_UM12_17_line4, M12_UM12_17_PT6_NotB);
inv M12_UM12_17_PT6_Xo3_2(M12_ContPar, M12_UM12_17_PT6_NotC);
and3 M12_UM12_17_PT6_Xo3_3(M12_UM12_17_PT6_NotA, M12_UM12_17_PT6_NotB, M12_ContPar, M12_UM12_17_PT6_line3);
and3 M12_UM12_17_PT6_Xo3_4(M12_UM12_17_PT6_NotA, M12_UM12_17_line4, M12_UM12_17_PT6_NotC, M12_UM12_17_PT6_line4);
and3 M12_UM12_17_PT6_Xo3_5(M12_UM12_17_line3, M12_UM12_17_PT6_NotB, M12_UM12_17_PT6_NotC, M12_UM12_17_PT6_line5);
and3 M12_UM12_17_PT6_Xo3_6(M12_UM12_17_line3, M12_UM12_17_line4, M12_ContPar, M12_UM12_17_PT6_line6);
nor2 M12_UM12_17_PT6_Xo3_7(M12_UM12_17_PT6_line3, M12_UM12_17_PT6_line4, M12_UM12_17_PT6_line7);
nor2 M12_UM12_17_PT6_Xo3_8(M12_UM12_17_PT6_line5, M12_UM12_17_PT6_line6, M12_UM12_17_PT6_line8);
nand2 M12_UM12_17_PT6_Xo3_9(M12_UM12_17_PT6_line7, M12_UM12_17_PT6_line8, M12_UM12_17_line6);
inv M12_UM12_17_PT7_Xo0(M12_UM12_17_line5, M12_UM12_17_PT7_NotA);
inv M12_UM12_17_PT7_Xo1(M12_UM12_17_line6, M12_UM12_17_PT7_NotB);
nand2 M12_UM12_17_PT7_Xo2(M12_UM12_17_PT7_NotA, M12_UM12_17_line6, M12_UM12_17_PT7_line2);
nand2 M12_UM12_17_PT7_Xo3(M12_UM12_17_PT7_NotB, M12_UM12_17_line5, M12_UM12_17_PT7_line3);
nand2 M12_UM12_17_PT7_Xo4(M12_UM12_17_PT7_line2, M12_UM12_17_PT7_line3, M12_EvenParZ_Cont);
inv M12_UM12_18(M12_EvenParA, out351);
inv M12_UM12_19(M12_EvenParB, out358);
inv M12_UM12_20(M12_EvenParZ, out402);
inv M12_UM12_21(M12_EvenParZ_Cont, out405);
inv M13_UM13_0_Inv8_0_Inv4_0(in116, M13_Not_Abus_0);
inv M13_UM13_0_Inv8_0_Inv4_1(in107, M13_Not_Abus_1);
inv M13_UM13_0_Inv8_0_Inv4_2(in97, M13_Not_Abus_2);
inv M13_UM13_0_Inv8_0_Inv4_3(in87, M13_Not_Abus_3);
inv M13_UM13_0_Inv8_1_Inv4_0(in77, M13_Not_Abus_4);
inv M13_UM13_0_Inv8_1_Inv4_1(in68, M13_Not_Abus_5);
inv M13_UM13_0_Inv8_1_Inv4_2(in58, M13_Not_Abus_6);
inv M13_UM13_0_Inv8_1_Inv4_3(in50, M13_Not_Abus_7);
inv M13_UM13_1_Xo0(in68, M13_UM13_1_NotA);
inv M13_UM13_1_Xo1(in58, M13_UM13_1_NotB);
nand2 M13_UM13_1_Xo2(M13_UM13_1_NotA, in58, M13_UM13_1_line2);
nand2 M13_UM13_1_Xo3(M13_UM13_1_NotB, in68, M13_UM13_1_line3);
nand2 M13_UM13_1_Xo4(M13_UM13_1_line2, M13_UM13_1_line3, M13_tmp0);
and3 M13_UM13_2(M13_tmp0, in77, in50, M13_tmp1);
and2 M13_UM13_3(in68, M13_Not_Abus_7, M13_tmp2);
or2 M13_UM13_4(M13_tmp1, M13_tmp2, M13_Misc0_0);
inv M13_UM13_5_Xo0(in107, M13_UM13_5_NotA);
inv M13_UM13_5_Xo1(in97, M13_UM13_5_NotB);
nand2 M13_UM13_5_Xo2(M13_UM13_5_NotA, in97, M13_UM13_5_line2);
nand2 M13_UM13_5_Xo3(M13_UM13_5_NotB, in107, M13_UM13_5_line3);
nand2 M13_UM13_5_Xo4(M13_UM13_5_line2, M13_UM13_5_line3, M13_tmp3);
and2 M13_UM13_6(in116, M13_tmp3, M13_Misc0_1);
inv M13_UM13_7(in13, M13_NotCont1);
inv M13_UM13_8(in41, M13_NotCont5);
nand2 M13_UM13_9(in1, M13_NotCont1, M13_ContHi_Misc0);
nand3 M13_UM13_10(in1, in13, in20, M13_ContLo_Misc0);
inv M13_UM13_11_Mux3c_0(M13_ContHi_Misc0, M13_UM13_11_NotContHi);
inv M13_UM13_11_Mux3c_1(M13_ContLo_Misc0, M13_UM13_11_NotContLo);
and2 M13_UM13_11_Mux3c_2(M13_Misc0_0, M13_UM13_11_NotContHi, M13_UM13_11_line2);
and2 M13_UM13_11_Mux3c_3(M13_Misc0_1, M13_UM13_11_NotContLo, M13_UM13_11_line3);
and2 M13_UM13_11_Mux3c_4(M13_ContHi_Misc0, M13_ContLo_Misc0, M13_UM13_11_line4);
and2 M13_UM13_11_Mux3c_5(M13_UM13_11_line4, Overflow, M13_UM13_11_line5);
or3 M13_UM13_11_Mux3c_6(M13_UM13_11_line2, M13_UM13_11_line3, M13_UM13_11_line5, out367);
or2 M13_UM13_12(in68, in58, M13_tmp4);
and2 M13_UM13_13(in50, M13_tmp4, M13_Misc1_0);
and4 M13_UM13_14(M13_Not_Abus_0, M13_Not_Abus_1, M13_Not_Abus_2, M13_Not_Abus_3, M13_Misc1_2);
nand4 M13_UM13_27(in1, M13_NotCont1, in20, M13_NotCont5, M13_ContHi_Misc1);
inv M13_UM13_28_Mux3c_0(M13_ContHi_Misc1, M13_UM13_28_NotContHi);
inv M13_UM13_28_Mux3c_1(in1, M13_UM13_28_NotContLo);
and2 M13_UM13_28_Mux3c_2(M13_Misc1_0, M13_UM13_28_NotContHi, M13_UM13_28_line2);
and2 M13_UM13_28_Mux3c_3(Carry4, M13_UM13_28_NotContLo, M13_UM13_28_line3);
and2 M13_UM13_28_Mux3c_4(M13_ContHi_Misc1, in1, M13_UM13_28_line4);
and2 M13_UM13_28_Mux3c_5(M13_UM13_28_line4, M13_Misc1_2, M13_UM13_28_line5);
or3 M13_UM13_28_Mux3c_6(M13_UM13_28_line2, M13_UM13_28_line3, M13_UM13_28_line5, out364);
or2 M13_UM13_29(in264, in257, M13_tmp5);
and2 M13_UM13_30(in250, M13_tmp5, M13_Misc2_1);
nand2 M13_UM13_31(in116, in270, M13_pr0);
nand2 M13_UM13_32(in107, in264, M13_pr1);
nand2 M13_UM13_33(in97, in257, M13_pr2);
nand2 M13_UM13_34(in87, in250, M13_pr3);
nand2 M13_UM13_35(in77, in244, M13_pr4);
nand2 M13_UM13_36(in68, in238, M13_pr5);
nand2 M13_UM13_37(in58, in232, M13_pr6);
nand2 M13_UM13_38(in50, in226, M13_pr7);
and4 M13_UM13_39(M13_pr0, M13_pr1, M13_pr2, M13_pr3, M13_pr3_0);
and4 M13_UM13_40(M13_pr4, M13_pr5, M13_pr6, M13_pr7, M13_pr7_4);
nand2 M13_UM13_41(M13_pr3_0, M13_pr7_4, M13_Misc2_2);
nand3 M13_UM13_42(in1, M13_NotCont1, in20, M13_ContLo_Misc2);
inv M13_UM13_43_Mux3c_0(M13_ContLo_Misc0, M13_UM13_43_NotContHi);
inv M13_UM13_43_Mux3c_1(M13_ContLo_Misc2, M13_UM13_43_NotContLo);
and2 M13_UM13_43_Mux3c_2(M13_Misc1_0, M13_UM13_43_NotContHi, M13_UM13_43_line2);
and2 M13_UM13_43_Mux3c_3(M13_Misc2_1, M13_UM13_43_NotContLo, M13_UM13_43_line3);
and2 M13_UM13_43_Mux3c_4(M13_ContLo_Misc0, M13_ContLo_Misc2, M13_UM13_43_line4);
and2 M13_UM13_43_Mux3c_5(M13_UM13_43_line4, M13_Misc2_2, M13_UM13_43_line5);
or3 M13_UM13_43_Mux3c_6(M13_UM13_43_line2, M13_UM13_43_line3, M13_UM13_43_line5, M13_NotMiscOuts2);
inv M13_UM13_43_1(M13_NotMiscOuts2, out361);
or2 M13_UM13_44(in107, in97, M13_tmp6);
and2 M13_UM13_45(in87, M13_tmp6, M13_tmp7);
inv M13_UM13_46(M13_tmp7, out355);
and4 M13_UM13_47(M13_Not_Abus_4, M13_Not_Abus_5, M13_Not_Abus_6, M13_Not_Abus_7, out353);

assign out399 = XCarrybus_2;
assign gnd = 1'b0;

endmodule
